
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MAC_32x16_8 IS
PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7, input_row_8, input_row_9, 
	input_row_10, input_row_11, input_row_12, input_row_13, input_row_14, input_row_15, input_row_16, input_row_17, input_row_18, input_row_19, 
	input_row_20, input_row_21, input_row_22, input_row_23, input_row_24, input_row_25, input_row_26, input_row_27, input_row_28, input_row_29, 
	input_row_30, input_row_31: IN STD_LOGIC_VECTOR(7 downto 0);
	input_col_0, input_col_1, input_col_2, input_col_3, input_col_4, input_col_5, input_col_6, input_col_7, input_col_8, input_col_9, 
	input_col_10, input_col_11, input_col_12, input_col_13, input_col_14, input_col_15: IN STD_LOGIC_VECTOR(7 downto 0);
	SEL_mux: IN STD_LOGIC_VECTOR(3 downto 0);
	CLK, RST_n, ENABLE : IN STD_LOGIC;
	output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7, output_row_8, output_row_9, 
	output_row_10, output_row_11, output_row_12, output_row_13, output_row_14, output_row_15, output_row_16, output_row_17, output_row_18, output_row_19, 
	output_row_20, output_row_21, output_row_22, output_row_23, output_row_24, output_row_25, output_row_26, output_row_27, output_row_28, output_row_29, 
	output_row_30, output_row_31: OUT STD_LOGIC_VECTOR(31 downto 0)
);
END MAC_32x16_8;

ARCHITECTURE behaviour OF  MAC_32x16_8 IS

	COMPONENT MAC IS
	GENERIC (data_size : POSITIVE := 2;
	 acc_size : POSITIVE := 16 );
	PORT( data_in_A, data_in_B  : IN STD_LOGIC_VECTOR(data_size-1 downto 0);
		CLK, RST_n, ENABLE 	: IN STD_LOGIC;
		data_out    			: OUT STD_LOGIC_VECTOR(acc_size-1 downto 0));
	END COMPONENT;

	COMPONENT mux_16to1_nbit IS
	GENERIC ( N : POSITIVE :=2);
	PORT(
		I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, 
		I10, I11, I12, I13, I14, I15: IN STD_LOGIC_VECTOR(N-1 downto 0);
		SEL_mux  : IN STD_LOGIC_VECTOR(3 downto 0);
		O    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
	END COMPONENT;


	SIGNAL output_MAC_0_0, output_MAC_0_1, output_MAC_0_2, output_MAC_0_3, output_MAC_0_4, output_MAC_0_5, output_MAC_0_6, output_MAC_0_7, output_MAC_0_8, output_MAC_0_9, 
		output_MAC_0_10, output_MAC_0_11, output_MAC_0_12, output_MAC_0_13, output_MAC_0_14, output_MAC_0_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_1_0, output_MAC_1_1, output_MAC_1_2, output_MAC_1_3, output_MAC_1_4, output_MAC_1_5, output_MAC_1_6, output_MAC_1_7, output_MAC_1_8, output_MAC_1_9, 
		output_MAC_1_10, output_MAC_1_11, output_MAC_1_12, output_MAC_1_13, output_MAC_1_14, output_MAC_1_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_2_0, output_MAC_2_1, output_MAC_2_2, output_MAC_2_3, output_MAC_2_4, output_MAC_2_5, output_MAC_2_6, output_MAC_2_7, output_MAC_2_8, output_MAC_2_9, 
		output_MAC_2_10, output_MAC_2_11, output_MAC_2_12, output_MAC_2_13, output_MAC_2_14, output_MAC_2_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_3_0, output_MAC_3_1, output_MAC_3_2, output_MAC_3_3, output_MAC_3_4, output_MAC_3_5, output_MAC_3_6, output_MAC_3_7, output_MAC_3_8, output_MAC_3_9, 
		output_MAC_3_10, output_MAC_3_11, output_MAC_3_12, output_MAC_3_13, output_MAC_3_14, output_MAC_3_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_4_0, output_MAC_4_1, output_MAC_4_2, output_MAC_4_3, output_MAC_4_4, output_MAC_4_5, output_MAC_4_6, output_MAC_4_7, output_MAC_4_8, output_MAC_4_9, 
		output_MAC_4_10, output_MAC_4_11, output_MAC_4_12, output_MAC_4_13, output_MAC_4_14, output_MAC_4_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_5_0, output_MAC_5_1, output_MAC_5_2, output_MAC_5_3, output_MAC_5_4, output_MAC_5_5, output_MAC_5_6, output_MAC_5_7, output_MAC_5_8, output_MAC_5_9, 
		output_MAC_5_10, output_MAC_5_11, output_MAC_5_12, output_MAC_5_13, output_MAC_5_14, output_MAC_5_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_6_0, output_MAC_6_1, output_MAC_6_2, output_MAC_6_3, output_MAC_6_4, output_MAC_6_5, output_MAC_6_6, output_MAC_6_7, output_MAC_6_8, output_MAC_6_9, 
		output_MAC_6_10, output_MAC_6_11, output_MAC_6_12, output_MAC_6_13, output_MAC_6_14, output_MAC_6_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_7_0, output_MAC_7_1, output_MAC_7_2, output_MAC_7_3, output_MAC_7_4, output_MAC_7_5, output_MAC_7_6, output_MAC_7_7, output_MAC_7_8, output_MAC_7_9, 
		output_MAC_7_10, output_MAC_7_11, output_MAC_7_12, output_MAC_7_13, output_MAC_7_14, output_MAC_7_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_8_0, output_MAC_8_1, output_MAC_8_2, output_MAC_8_3, output_MAC_8_4, output_MAC_8_5, output_MAC_8_6, output_MAC_8_7, output_MAC_8_8, output_MAC_8_9, 
		output_MAC_8_10, output_MAC_8_11, output_MAC_8_12, output_MAC_8_13, output_MAC_8_14, output_MAC_8_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_9_0, output_MAC_9_1, output_MAC_9_2, output_MAC_9_3, output_MAC_9_4, output_MAC_9_5, output_MAC_9_6, output_MAC_9_7, output_MAC_9_8, output_MAC_9_9, 
		output_MAC_9_10, output_MAC_9_11, output_MAC_9_12, output_MAC_9_13, output_MAC_9_14, output_MAC_9_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_10_0, output_MAC_10_1, output_MAC_10_2, output_MAC_10_3, output_MAC_10_4, output_MAC_10_5, output_MAC_10_6, output_MAC_10_7, output_MAC_10_8, output_MAC_10_9, 
		output_MAC_10_10, output_MAC_10_11, output_MAC_10_12, output_MAC_10_13, output_MAC_10_14, output_MAC_10_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_11_0, output_MAC_11_1, output_MAC_11_2, output_MAC_11_3, output_MAC_11_4, output_MAC_11_5, output_MAC_11_6, output_MAC_11_7, output_MAC_11_8, output_MAC_11_9, 
		output_MAC_11_10, output_MAC_11_11, output_MAC_11_12, output_MAC_11_13, output_MAC_11_14, output_MAC_11_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_12_0, output_MAC_12_1, output_MAC_12_2, output_MAC_12_3, output_MAC_12_4, output_MAC_12_5, output_MAC_12_6, output_MAC_12_7, output_MAC_12_8, output_MAC_12_9, 
		output_MAC_12_10, output_MAC_12_11, output_MAC_12_12, output_MAC_12_13, output_MAC_12_14, output_MAC_12_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_13_0, output_MAC_13_1, output_MAC_13_2, output_MAC_13_3, output_MAC_13_4, output_MAC_13_5, output_MAC_13_6, output_MAC_13_7, output_MAC_13_8, output_MAC_13_9, 
		output_MAC_13_10, output_MAC_13_11, output_MAC_13_12, output_MAC_13_13, output_MAC_13_14, output_MAC_13_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_14_0, output_MAC_14_1, output_MAC_14_2, output_MAC_14_3, output_MAC_14_4, output_MAC_14_5, output_MAC_14_6, output_MAC_14_7, output_MAC_14_8, output_MAC_14_9, 
		output_MAC_14_10, output_MAC_14_11, output_MAC_14_12, output_MAC_14_13, output_MAC_14_14, output_MAC_14_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_15_0, output_MAC_15_1, output_MAC_15_2, output_MAC_15_3, output_MAC_15_4, output_MAC_15_5, output_MAC_15_6, output_MAC_15_7, output_MAC_15_8, output_MAC_15_9, 
		output_MAC_15_10, output_MAC_15_11, output_MAC_15_12, output_MAC_15_13, output_MAC_15_14, output_MAC_15_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_16_0, output_MAC_16_1, output_MAC_16_2, output_MAC_16_3, output_MAC_16_4, output_MAC_16_5, output_MAC_16_6, output_MAC_16_7, output_MAC_16_8, output_MAC_16_9, 
		output_MAC_16_10, output_MAC_16_11, output_MAC_16_12, output_MAC_16_13, output_MAC_16_14, output_MAC_16_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_17_0, output_MAC_17_1, output_MAC_17_2, output_MAC_17_3, output_MAC_17_4, output_MAC_17_5, output_MAC_17_6, output_MAC_17_7, output_MAC_17_8, output_MAC_17_9, 
		output_MAC_17_10, output_MAC_17_11, output_MAC_17_12, output_MAC_17_13, output_MAC_17_14, output_MAC_17_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_18_0, output_MAC_18_1, output_MAC_18_2, output_MAC_18_3, output_MAC_18_4, output_MAC_18_5, output_MAC_18_6, output_MAC_18_7, output_MAC_18_8, output_MAC_18_9, 
		output_MAC_18_10, output_MAC_18_11, output_MAC_18_12, output_MAC_18_13, output_MAC_18_14, output_MAC_18_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_19_0, output_MAC_19_1, output_MAC_19_2, output_MAC_19_3, output_MAC_19_4, output_MAC_19_5, output_MAC_19_6, output_MAC_19_7, output_MAC_19_8, output_MAC_19_9, 
		output_MAC_19_10, output_MAC_19_11, output_MAC_19_12, output_MAC_19_13, output_MAC_19_14, output_MAC_19_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_20_0, output_MAC_20_1, output_MAC_20_2, output_MAC_20_3, output_MAC_20_4, output_MAC_20_5, output_MAC_20_6, output_MAC_20_7, output_MAC_20_8, output_MAC_20_9, 
		output_MAC_20_10, output_MAC_20_11, output_MAC_20_12, output_MAC_20_13, output_MAC_20_14, output_MAC_20_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_21_0, output_MAC_21_1, output_MAC_21_2, output_MAC_21_3, output_MAC_21_4, output_MAC_21_5, output_MAC_21_6, output_MAC_21_7, output_MAC_21_8, output_MAC_21_9, 
		output_MAC_21_10, output_MAC_21_11, output_MAC_21_12, output_MAC_21_13, output_MAC_21_14, output_MAC_21_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_22_0, output_MAC_22_1, output_MAC_22_2, output_MAC_22_3, output_MAC_22_4, output_MAC_22_5, output_MAC_22_6, output_MAC_22_7, output_MAC_22_8, output_MAC_22_9, 
		output_MAC_22_10, output_MAC_22_11, output_MAC_22_12, output_MAC_22_13, output_MAC_22_14, output_MAC_22_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_23_0, output_MAC_23_1, output_MAC_23_2, output_MAC_23_3, output_MAC_23_4, output_MAC_23_5, output_MAC_23_6, output_MAC_23_7, output_MAC_23_8, output_MAC_23_9, 
		output_MAC_23_10, output_MAC_23_11, output_MAC_23_12, output_MAC_23_13, output_MAC_23_14, output_MAC_23_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_24_0, output_MAC_24_1, output_MAC_24_2, output_MAC_24_3, output_MAC_24_4, output_MAC_24_5, output_MAC_24_6, output_MAC_24_7, output_MAC_24_8, output_MAC_24_9, 
		output_MAC_24_10, output_MAC_24_11, output_MAC_24_12, output_MAC_24_13, output_MAC_24_14, output_MAC_24_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_25_0, output_MAC_25_1, output_MAC_25_2, output_MAC_25_3, output_MAC_25_4, output_MAC_25_5, output_MAC_25_6, output_MAC_25_7, output_MAC_25_8, output_MAC_25_9, 
		output_MAC_25_10, output_MAC_25_11, output_MAC_25_12, output_MAC_25_13, output_MAC_25_14, output_MAC_25_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_26_0, output_MAC_26_1, output_MAC_26_2, output_MAC_26_3, output_MAC_26_4, output_MAC_26_5, output_MAC_26_6, output_MAC_26_7, output_MAC_26_8, output_MAC_26_9, 
		output_MAC_26_10, output_MAC_26_11, output_MAC_26_12, output_MAC_26_13, output_MAC_26_14, output_MAC_26_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_27_0, output_MAC_27_1, output_MAC_27_2, output_MAC_27_3, output_MAC_27_4, output_MAC_27_5, output_MAC_27_6, output_MAC_27_7, output_MAC_27_8, output_MAC_27_9, 
		output_MAC_27_10, output_MAC_27_11, output_MAC_27_12, output_MAC_27_13, output_MAC_27_14, output_MAC_27_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_28_0, output_MAC_28_1, output_MAC_28_2, output_MAC_28_3, output_MAC_28_4, output_MAC_28_5, output_MAC_28_6, output_MAC_28_7, output_MAC_28_8, output_MAC_28_9, 
		output_MAC_28_10, output_MAC_28_11, output_MAC_28_12, output_MAC_28_13, output_MAC_28_14, output_MAC_28_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_29_0, output_MAC_29_1, output_MAC_29_2, output_MAC_29_3, output_MAC_29_4, output_MAC_29_5, output_MAC_29_6, output_MAC_29_7, output_MAC_29_8, output_MAC_29_9, 
		output_MAC_29_10, output_MAC_29_11, output_MAC_29_12, output_MAC_29_13, output_MAC_29_14, output_MAC_29_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_30_0, output_MAC_30_1, output_MAC_30_2, output_MAC_30_3, output_MAC_30_4, output_MAC_30_5, output_MAC_30_6, output_MAC_30_7, output_MAC_30_8, output_MAC_30_9, 
		output_MAC_30_10, output_MAC_30_11, output_MAC_30_12, output_MAC_30_13, output_MAC_30_14, output_MAC_30_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_31_0, output_MAC_31_1, output_MAC_31_2, output_MAC_31_3, output_MAC_31_4, output_MAC_31_5, output_MAC_31_6, output_MAC_31_7, output_MAC_31_8, output_MAC_31_9, 
		output_MAC_31_10, output_MAC_31_11, output_MAC_31_12, output_MAC_31_13, output_MAC_31_14, output_MAC_31_15: STD_LOGIC_VECTOR(31 downto 0);

BEGIN

	MAC_0_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_0, data_out=>output_MAC_0_0);
	MAC_0_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_1, data_out=>output_MAC_0_1);
	MAC_0_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_2, data_out=>output_MAC_0_2);
	MAC_0_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_3, data_out=>output_MAC_0_3);
	MAC_0_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_4, data_out=>output_MAC_0_4);
	MAC_0_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_5, data_out=>output_MAC_0_5);
	MAC_0_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_6, data_out=>output_MAC_0_6);
	MAC_0_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_7, data_out=>output_MAC_0_7);
	MAC_0_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_8, data_out=>output_MAC_0_8);
	MAC_0_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_9, data_out=>output_MAC_0_9);
	MAC_0_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_10, data_out=>output_MAC_0_10);
	MAC_0_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_11, data_out=>output_MAC_0_11);
	MAC_0_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_12, data_out=>output_MAC_0_12);
	MAC_0_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_13, data_out=>output_MAC_0_13);
	MAC_0_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_14, data_out=>output_MAC_0_14);
	MAC_0_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_15, data_out=>output_MAC_0_15);
	MAC_1_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_0, data_out=>output_MAC_1_0);
	MAC_1_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_1, data_out=>output_MAC_1_1);
	MAC_1_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_2, data_out=>output_MAC_1_2);
	MAC_1_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_3, data_out=>output_MAC_1_3);
	MAC_1_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_4, data_out=>output_MAC_1_4);
	MAC_1_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_5, data_out=>output_MAC_1_5);
	MAC_1_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_6, data_out=>output_MAC_1_6);
	MAC_1_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_7, data_out=>output_MAC_1_7);
	MAC_1_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_8, data_out=>output_MAC_1_8);
	MAC_1_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_9, data_out=>output_MAC_1_9);
	MAC_1_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_10, data_out=>output_MAC_1_10);
	MAC_1_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_11, data_out=>output_MAC_1_11);
	MAC_1_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_12, data_out=>output_MAC_1_12);
	MAC_1_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_13, data_out=>output_MAC_1_13);
	MAC_1_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_14, data_out=>output_MAC_1_14);
	MAC_1_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_15, data_out=>output_MAC_1_15);
	MAC_2_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_0, data_out=>output_MAC_2_0);
	MAC_2_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_1, data_out=>output_MAC_2_1);
	MAC_2_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_2, data_out=>output_MAC_2_2);
	MAC_2_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_3, data_out=>output_MAC_2_3);
	MAC_2_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_4, data_out=>output_MAC_2_4);
	MAC_2_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_5, data_out=>output_MAC_2_5);
	MAC_2_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_6, data_out=>output_MAC_2_6);
	MAC_2_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_7, data_out=>output_MAC_2_7);
	MAC_2_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_8, data_out=>output_MAC_2_8);
	MAC_2_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_9, data_out=>output_MAC_2_9);
	MAC_2_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_10, data_out=>output_MAC_2_10);
	MAC_2_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_11, data_out=>output_MAC_2_11);
	MAC_2_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_12, data_out=>output_MAC_2_12);
	MAC_2_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_13, data_out=>output_MAC_2_13);
	MAC_2_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_14, data_out=>output_MAC_2_14);
	MAC_2_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_15, data_out=>output_MAC_2_15);
	MAC_3_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_0, data_out=>output_MAC_3_0);
	MAC_3_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_1, data_out=>output_MAC_3_1);
	MAC_3_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_2, data_out=>output_MAC_3_2);
	MAC_3_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_3, data_out=>output_MAC_3_3);
	MAC_3_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_4, data_out=>output_MAC_3_4);
	MAC_3_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_5, data_out=>output_MAC_3_5);
	MAC_3_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_6, data_out=>output_MAC_3_6);
	MAC_3_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_7, data_out=>output_MAC_3_7);
	MAC_3_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_8, data_out=>output_MAC_3_8);
	MAC_3_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_9, data_out=>output_MAC_3_9);
	MAC_3_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_10, data_out=>output_MAC_3_10);
	MAC_3_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_11, data_out=>output_MAC_3_11);
	MAC_3_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_12, data_out=>output_MAC_3_12);
	MAC_3_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_13, data_out=>output_MAC_3_13);
	MAC_3_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_14, data_out=>output_MAC_3_14);
	MAC_3_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_15, data_out=>output_MAC_3_15);
	MAC_4_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_0, data_out=>output_MAC_4_0);
	MAC_4_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_1, data_out=>output_MAC_4_1);
	MAC_4_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_2, data_out=>output_MAC_4_2);
	MAC_4_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_3, data_out=>output_MAC_4_3);
	MAC_4_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_4, data_out=>output_MAC_4_4);
	MAC_4_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_5, data_out=>output_MAC_4_5);
	MAC_4_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_6, data_out=>output_MAC_4_6);
	MAC_4_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_7, data_out=>output_MAC_4_7);
	MAC_4_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_8, data_out=>output_MAC_4_8);
	MAC_4_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_9, data_out=>output_MAC_4_9);
	MAC_4_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_10, data_out=>output_MAC_4_10);
	MAC_4_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_11, data_out=>output_MAC_4_11);
	MAC_4_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_12, data_out=>output_MAC_4_12);
	MAC_4_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_13, data_out=>output_MAC_4_13);
	MAC_4_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_14, data_out=>output_MAC_4_14);
	MAC_4_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_15, data_out=>output_MAC_4_15);
	MAC_5_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_0, data_out=>output_MAC_5_0);
	MAC_5_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_1, data_out=>output_MAC_5_1);
	MAC_5_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_2, data_out=>output_MAC_5_2);
	MAC_5_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_3, data_out=>output_MAC_5_3);
	MAC_5_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_4, data_out=>output_MAC_5_4);
	MAC_5_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_5, data_out=>output_MAC_5_5);
	MAC_5_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_6, data_out=>output_MAC_5_6);
	MAC_5_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_7, data_out=>output_MAC_5_7);
	MAC_5_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_8, data_out=>output_MAC_5_8);
	MAC_5_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_9, data_out=>output_MAC_5_9);
	MAC_5_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_10, data_out=>output_MAC_5_10);
	MAC_5_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_11, data_out=>output_MAC_5_11);
	MAC_5_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_12, data_out=>output_MAC_5_12);
	MAC_5_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_13, data_out=>output_MAC_5_13);
	MAC_5_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_14, data_out=>output_MAC_5_14);
	MAC_5_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_15, data_out=>output_MAC_5_15);
	MAC_6_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_0, data_out=>output_MAC_6_0);
	MAC_6_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_1, data_out=>output_MAC_6_1);
	MAC_6_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_2, data_out=>output_MAC_6_2);
	MAC_6_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_3, data_out=>output_MAC_6_3);
	MAC_6_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_4, data_out=>output_MAC_6_4);
	MAC_6_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_5, data_out=>output_MAC_6_5);
	MAC_6_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_6, data_out=>output_MAC_6_6);
	MAC_6_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_7, data_out=>output_MAC_6_7);
	MAC_6_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_8, data_out=>output_MAC_6_8);
	MAC_6_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_9, data_out=>output_MAC_6_9);
	MAC_6_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_10, data_out=>output_MAC_6_10);
	MAC_6_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_11, data_out=>output_MAC_6_11);
	MAC_6_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_12, data_out=>output_MAC_6_12);
	MAC_6_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_13, data_out=>output_MAC_6_13);
	MAC_6_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_14, data_out=>output_MAC_6_14);
	MAC_6_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_15, data_out=>output_MAC_6_15);
	MAC_7_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_0, data_out=>output_MAC_7_0);
	MAC_7_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_1, data_out=>output_MAC_7_1);
	MAC_7_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_2, data_out=>output_MAC_7_2);
	MAC_7_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_3, data_out=>output_MAC_7_3);
	MAC_7_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_4, data_out=>output_MAC_7_4);
	MAC_7_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_5, data_out=>output_MAC_7_5);
	MAC_7_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_6, data_out=>output_MAC_7_6);
	MAC_7_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_7, data_out=>output_MAC_7_7);
	MAC_7_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_8, data_out=>output_MAC_7_8);
	MAC_7_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_9, data_out=>output_MAC_7_9);
	MAC_7_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_10, data_out=>output_MAC_7_10);
	MAC_7_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_11, data_out=>output_MAC_7_11);
	MAC_7_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_12, data_out=>output_MAC_7_12);
	MAC_7_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_13, data_out=>output_MAC_7_13);
	MAC_7_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_14, data_out=>output_MAC_7_14);
	MAC_7_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_15, data_out=>output_MAC_7_15);
	MAC_8_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_0, data_out=>output_MAC_8_0);
	MAC_8_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_1, data_out=>output_MAC_8_1);
	MAC_8_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_2, data_out=>output_MAC_8_2);
	MAC_8_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_3, data_out=>output_MAC_8_3);
	MAC_8_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_4, data_out=>output_MAC_8_4);
	MAC_8_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_5, data_out=>output_MAC_8_5);
	MAC_8_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_6, data_out=>output_MAC_8_6);
	MAC_8_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_7, data_out=>output_MAC_8_7);
	MAC_8_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_8, data_out=>output_MAC_8_8);
	MAC_8_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_9, data_out=>output_MAC_8_9);
	MAC_8_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_10, data_out=>output_MAC_8_10);
	MAC_8_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_11, data_out=>output_MAC_8_11);
	MAC_8_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_12, data_out=>output_MAC_8_12);
	MAC_8_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_13, data_out=>output_MAC_8_13);
	MAC_8_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_14, data_out=>output_MAC_8_14);
	MAC_8_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_15, data_out=>output_MAC_8_15);
	MAC_9_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_0, data_out=>output_MAC_9_0);
	MAC_9_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_1, data_out=>output_MAC_9_1);
	MAC_9_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_2, data_out=>output_MAC_9_2);
	MAC_9_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_3, data_out=>output_MAC_9_3);
	MAC_9_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_4, data_out=>output_MAC_9_4);
	MAC_9_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_5, data_out=>output_MAC_9_5);
	MAC_9_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_6, data_out=>output_MAC_9_6);
	MAC_9_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_7, data_out=>output_MAC_9_7);
	MAC_9_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_8, data_out=>output_MAC_9_8);
	MAC_9_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_9, data_out=>output_MAC_9_9);
	MAC_9_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_10, data_out=>output_MAC_9_10);
	MAC_9_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_11, data_out=>output_MAC_9_11);
	MAC_9_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_12, data_out=>output_MAC_9_12);
	MAC_9_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_13, data_out=>output_MAC_9_13);
	MAC_9_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_14, data_out=>output_MAC_9_14);
	MAC_9_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_15, data_out=>output_MAC_9_15);
	MAC_10_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_0, data_out=>output_MAC_10_0);
	MAC_10_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_1, data_out=>output_MAC_10_1);
	MAC_10_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_2, data_out=>output_MAC_10_2);
	MAC_10_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_3, data_out=>output_MAC_10_3);
	MAC_10_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_4, data_out=>output_MAC_10_4);
	MAC_10_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_5, data_out=>output_MAC_10_5);
	MAC_10_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_6, data_out=>output_MAC_10_6);
	MAC_10_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_7, data_out=>output_MAC_10_7);
	MAC_10_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_8, data_out=>output_MAC_10_8);
	MAC_10_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_9, data_out=>output_MAC_10_9);
	MAC_10_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_10, data_out=>output_MAC_10_10);
	MAC_10_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_11, data_out=>output_MAC_10_11);
	MAC_10_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_12, data_out=>output_MAC_10_12);
	MAC_10_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_13, data_out=>output_MAC_10_13);
	MAC_10_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_14, data_out=>output_MAC_10_14);
	MAC_10_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_15, data_out=>output_MAC_10_15);
	MAC_11_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_0, data_out=>output_MAC_11_0);
	MAC_11_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_1, data_out=>output_MAC_11_1);
	MAC_11_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_2, data_out=>output_MAC_11_2);
	MAC_11_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_3, data_out=>output_MAC_11_3);
	MAC_11_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_4, data_out=>output_MAC_11_4);
	MAC_11_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_5, data_out=>output_MAC_11_5);
	MAC_11_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_6, data_out=>output_MAC_11_6);
	MAC_11_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_7, data_out=>output_MAC_11_7);
	MAC_11_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_8, data_out=>output_MAC_11_8);
	MAC_11_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_9, data_out=>output_MAC_11_9);
	MAC_11_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_10, data_out=>output_MAC_11_10);
	MAC_11_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_11, data_out=>output_MAC_11_11);
	MAC_11_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_12, data_out=>output_MAC_11_12);
	MAC_11_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_13, data_out=>output_MAC_11_13);
	MAC_11_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_14, data_out=>output_MAC_11_14);
	MAC_11_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_15, data_out=>output_MAC_11_15);
	MAC_12_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_0, data_out=>output_MAC_12_0);
	MAC_12_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_1, data_out=>output_MAC_12_1);
	MAC_12_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_2, data_out=>output_MAC_12_2);
	MAC_12_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_3, data_out=>output_MAC_12_3);
	MAC_12_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_4, data_out=>output_MAC_12_4);
	MAC_12_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_5, data_out=>output_MAC_12_5);
	MAC_12_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_6, data_out=>output_MAC_12_6);
	MAC_12_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_7, data_out=>output_MAC_12_7);
	MAC_12_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_8, data_out=>output_MAC_12_8);
	MAC_12_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_9, data_out=>output_MAC_12_9);
	MAC_12_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_10, data_out=>output_MAC_12_10);
	MAC_12_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_11, data_out=>output_MAC_12_11);
	MAC_12_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_12, data_out=>output_MAC_12_12);
	MAC_12_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_13, data_out=>output_MAC_12_13);
	MAC_12_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_14, data_out=>output_MAC_12_14);
	MAC_12_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_15, data_out=>output_MAC_12_15);
	MAC_13_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_0, data_out=>output_MAC_13_0);
	MAC_13_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_1, data_out=>output_MAC_13_1);
	MAC_13_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_2, data_out=>output_MAC_13_2);
	MAC_13_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_3, data_out=>output_MAC_13_3);
	MAC_13_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_4, data_out=>output_MAC_13_4);
	MAC_13_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_5, data_out=>output_MAC_13_5);
	MAC_13_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_6, data_out=>output_MAC_13_6);
	MAC_13_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_7, data_out=>output_MAC_13_7);
	MAC_13_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_8, data_out=>output_MAC_13_8);
	MAC_13_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_9, data_out=>output_MAC_13_9);
	MAC_13_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_10, data_out=>output_MAC_13_10);
	MAC_13_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_11, data_out=>output_MAC_13_11);
	MAC_13_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_12, data_out=>output_MAC_13_12);
	MAC_13_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_13, data_out=>output_MAC_13_13);
	MAC_13_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_14, data_out=>output_MAC_13_14);
	MAC_13_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_15, data_out=>output_MAC_13_15);
	MAC_14_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_0, data_out=>output_MAC_14_0);
	MAC_14_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_1, data_out=>output_MAC_14_1);
	MAC_14_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_2, data_out=>output_MAC_14_2);
	MAC_14_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_3, data_out=>output_MAC_14_3);
	MAC_14_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_4, data_out=>output_MAC_14_4);
	MAC_14_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_5, data_out=>output_MAC_14_5);
	MAC_14_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_6, data_out=>output_MAC_14_6);
	MAC_14_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_7, data_out=>output_MAC_14_7);
	MAC_14_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_8, data_out=>output_MAC_14_8);
	MAC_14_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_9, data_out=>output_MAC_14_9);
	MAC_14_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_10, data_out=>output_MAC_14_10);
	MAC_14_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_11, data_out=>output_MAC_14_11);
	MAC_14_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_12, data_out=>output_MAC_14_12);
	MAC_14_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_13, data_out=>output_MAC_14_13);
	MAC_14_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_14, data_out=>output_MAC_14_14);
	MAC_14_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_15, data_out=>output_MAC_14_15);
	MAC_15_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_0, data_out=>output_MAC_15_0);
	MAC_15_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_1, data_out=>output_MAC_15_1);
	MAC_15_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_2, data_out=>output_MAC_15_2);
	MAC_15_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_3, data_out=>output_MAC_15_3);
	MAC_15_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_4, data_out=>output_MAC_15_4);
	MAC_15_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_5, data_out=>output_MAC_15_5);
	MAC_15_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_6, data_out=>output_MAC_15_6);
	MAC_15_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_7, data_out=>output_MAC_15_7);
	MAC_15_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_8, data_out=>output_MAC_15_8);
	MAC_15_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_9, data_out=>output_MAC_15_9);
	MAC_15_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_10, data_out=>output_MAC_15_10);
	MAC_15_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_11, data_out=>output_MAC_15_11);
	MAC_15_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_12, data_out=>output_MAC_15_12);
	MAC_15_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_13, data_out=>output_MAC_15_13);
	MAC_15_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_14, data_out=>output_MAC_15_14);
	MAC_15_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_15, data_out=>output_MAC_15_15);
	MAC_16_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_0, data_out=>output_MAC_16_0);
	MAC_16_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_1, data_out=>output_MAC_16_1);
	MAC_16_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_2, data_out=>output_MAC_16_2);
	MAC_16_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_3, data_out=>output_MAC_16_3);
	MAC_16_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_4, data_out=>output_MAC_16_4);
	MAC_16_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_5, data_out=>output_MAC_16_5);
	MAC_16_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_6, data_out=>output_MAC_16_6);
	MAC_16_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_7, data_out=>output_MAC_16_7);
	MAC_16_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_8, data_out=>output_MAC_16_8);
	MAC_16_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_9, data_out=>output_MAC_16_9);
	MAC_16_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_10, data_out=>output_MAC_16_10);
	MAC_16_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_11, data_out=>output_MAC_16_11);
	MAC_16_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_12, data_out=>output_MAC_16_12);
	MAC_16_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_13, data_out=>output_MAC_16_13);
	MAC_16_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_14, data_out=>output_MAC_16_14);
	MAC_16_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_15, data_out=>output_MAC_16_15);
	MAC_17_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_0, data_out=>output_MAC_17_0);
	MAC_17_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_1, data_out=>output_MAC_17_1);
	MAC_17_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_2, data_out=>output_MAC_17_2);
	MAC_17_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_3, data_out=>output_MAC_17_3);
	MAC_17_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_4, data_out=>output_MAC_17_4);
	MAC_17_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_5, data_out=>output_MAC_17_5);
	MAC_17_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_6, data_out=>output_MAC_17_6);
	MAC_17_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_7, data_out=>output_MAC_17_7);
	MAC_17_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_8, data_out=>output_MAC_17_8);
	MAC_17_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_9, data_out=>output_MAC_17_9);
	MAC_17_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_10, data_out=>output_MAC_17_10);
	MAC_17_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_11, data_out=>output_MAC_17_11);
	MAC_17_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_12, data_out=>output_MAC_17_12);
	MAC_17_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_13, data_out=>output_MAC_17_13);
	MAC_17_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_14, data_out=>output_MAC_17_14);
	MAC_17_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_15, data_out=>output_MAC_17_15);
	MAC_18_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_0, data_out=>output_MAC_18_0);
	MAC_18_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_1, data_out=>output_MAC_18_1);
	MAC_18_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_2, data_out=>output_MAC_18_2);
	MAC_18_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_3, data_out=>output_MAC_18_3);
	MAC_18_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_4, data_out=>output_MAC_18_4);
	MAC_18_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_5, data_out=>output_MAC_18_5);
	MAC_18_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_6, data_out=>output_MAC_18_6);
	MAC_18_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_7, data_out=>output_MAC_18_7);
	MAC_18_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_8, data_out=>output_MAC_18_8);
	MAC_18_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_9, data_out=>output_MAC_18_9);
	MAC_18_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_10, data_out=>output_MAC_18_10);
	MAC_18_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_11, data_out=>output_MAC_18_11);
	MAC_18_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_12, data_out=>output_MAC_18_12);
	MAC_18_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_13, data_out=>output_MAC_18_13);
	MAC_18_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_14, data_out=>output_MAC_18_14);
	MAC_18_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_15, data_out=>output_MAC_18_15);
	MAC_19_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_0, data_out=>output_MAC_19_0);
	MAC_19_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_1, data_out=>output_MAC_19_1);
	MAC_19_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_2, data_out=>output_MAC_19_2);
	MAC_19_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_3, data_out=>output_MAC_19_3);
	MAC_19_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_4, data_out=>output_MAC_19_4);
	MAC_19_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_5, data_out=>output_MAC_19_5);
	MAC_19_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_6, data_out=>output_MAC_19_6);
	MAC_19_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_7, data_out=>output_MAC_19_7);
	MAC_19_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_8, data_out=>output_MAC_19_8);
	MAC_19_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_9, data_out=>output_MAC_19_9);
	MAC_19_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_10, data_out=>output_MAC_19_10);
	MAC_19_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_11, data_out=>output_MAC_19_11);
	MAC_19_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_12, data_out=>output_MAC_19_12);
	MAC_19_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_13, data_out=>output_MAC_19_13);
	MAC_19_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_14, data_out=>output_MAC_19_14);
	MAC_19_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_15, data_out=>output_MAC_19_15);
	MAC_20_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_0, data_out=>output_MAC_20_0);
	MAC_20_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_1, data_out=>output_MAC_20_1);
	MAC_20_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_2, data_out=>output_MAC_20_2);
	MAC_20_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_3, data_out=>output_MAC_20_3);
	MAC_20_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_4, data_out=>output_MAC_20_4);
	MAC_20_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_5, data_out=>output_MAC_20_5);
	MAC_20_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_6, data_out=>output_MAC_20_6);
	MAC_20_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_7, data_out=>output_MAC_20_7);
	MAC_20_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_8, data_out=>output_MAC_20_8);
	MAC_20_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_9, data_out=>output_MAC_20_9);
	MAC_20_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_10, data_out=>output_MAC_20_10);
	MAC_20_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_11, data_out=>output_MAC_20_11);
	MAC_20_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_12, data_out=>output_MAC_20_12);
	MAC_20_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_13, data_out=>output_MAC_20_13);
	MAC_20_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_14, data_out=>output_MAC_20_14);
	MAC_20_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_15, data_out=>output_MAC_20_15);
	MAC_21_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_0, data_out=>output_MAC_21_0);
	MAC_21_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_1, data_out=>output_MAC_21_1);
	MAC_21_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_2, data_out=>output_MAC_21_2);
	MAC_21_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_3, data_out=>output_MAC_21_3);
	MAC_21_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_4, data_out=>output_MAC_21_4);
	MAC_21_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_5, data_out=>output_MAC_21_5);
	MAC_21_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_6, data_out=>output_MAC_21_6);
	MAC_21_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_7, data_out=>output_MAC_21_7);
	MAC_21_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_8, data_out=>output_MAC_21_8);
	MAC_21_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_9, data_out=>output_MAC_21_9);
	MAC_21_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_10, data_out=>output_MAC_21_10);
	MAC_21_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_11, data_out=>output_MAC_21_11);
	MAC_21_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_12, data_out=>output_MAC_21_12);
	MAC_21_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_13, data_out=>output_MAC_21_13);
	MAC_21_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_14, data_out=>output_MAC_21_14);
	MAC_21_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_15, data_out=>output_MAC_21_15);
	MAC_22_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_0, data_out=>output_MAC_22_0);
	MAC_22_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_1, data_out=>output_MAC_22_1);
	MAC_22_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_2, data_out=>output_MAC_22_2);
	MAC_22_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_3, data_out=>output_MAC_22_3);
	MAC_22_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_4, data_out=>output_MAC_22_4);
	MAC_22_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_5, data_out=>output_MAC_22_5);
	MAC_22_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_6, data_out=>output_MAC_22_6);
	MAC_22_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_7, data_out=>output_MAC_22_7);
	MAC_22_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_8, data_out=>output_MAC_22_8);
	MAC_22_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_9, data_out=>output_MAC_22_9);
	MAC_22_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_10, data_out=>output_MAC_22_10);
	MAC_22_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_11, data_out=>output_MAC_22_11);
	MAC_22_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_12, data_out=>output_MAC_22_12);
	MAC_22_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_13, data_out=>output_MAC_22_13);
	MAC_22_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_14, data_out=>output_MAC_22_14);
	MAC_22_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_15, data_out=>output_MAC_22_15);
	MAC_23_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_0, data_out=>output_MAC_23_0);
	MAC_23_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_1, data_out=>output_MAC_23_1);
	MAC_23_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_2, data_out=>output_MAC_23_2);
	MAC_23_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_3, data_out=>output_MAC_23_3);
	MAC_23_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_4, data_out=>output_MAC_23_4);
	MAC_23_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_5, data_out=>output_MAC_23_5);
	MAC_23_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_6, data_out=>output_MAC_23_6);
	MAC_23_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_7, data_out=>output_MAC_23_7);
	MAC_23_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_8, data_out=>output_MAC_23_8);
	MAC_23_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_9, data_out=>output_MAC_23_9);
	MAC_23_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_10, data_out=>output_MAC_23_10);
	MAC_23_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_11, data_out=>output_MAC_23_11);
	MAC_23_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_12, data_out=>output_MAC_23_12);
	MAC_23_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_13, data_out=>output_MAC_23_13);
	MAC_23_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_14, data_out=>output_MAC_23_14);
	MAC_23_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_15, data_out=>output_MAC_23_15);
	MAC_24_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_0, data_out=>output_MAC_24_0);
	MAC_24_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_1, data_out=>output_MAC_24_1);
	MAC_24_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_2, data_out=>output_MAC_24_2);
	MAC_24_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_3, data_out=>output_MAC_24_3);
	MAC_24_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_4, data_out=>output_MAC_24_4);
	MAC_24_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_5, data_out=>output_MAC_24_5);
	MAC_24_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_6, data_out=>output_MAC_24_6);
	MAC_24_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_7, data_out=>output_MAC_24_7);
	MAC_24_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_8, data_out=>output_MAC_24_8);
	MAC_24_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_9, data_out=>output_MAC_24_9);
	MAC_24_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_10, data_out=>output_MAC_24_10);
	MAC_24_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_11, data_out=>output_MAC_24_11);
	MAC_24_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_12, data_out=>output_MAC_24_12);
	MAC_24_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_13, data_out=>output_MAC_24_13);
	MAC_24_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_14, data_out=>output_MAC_24_14);
	MAC_24_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_15, data_out=>output_MAC_24_15);
	MAC_25_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_0, data_out=>output_MAC_25_0);
	MAC_25_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_1, data_out=>output_MAC_25_1);
	MAC_25_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_2, data_out=>output_MAC_25_2);
	MAC_25_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_3, data_out=>output_MAC_25_3);
	MAC_25_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_4, data_out=>output_MAC_25_4);
	MAC_25_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_5, data_out=>output_MAC_25_5);
	MAC_25_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_6, data_out=>output_MAC_25_6);
	MAC_25_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_7, data_out=>output_MAC_25_7);
	MAC_25_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_8, data_out=>output_MAC_25_8);
	MAC_25_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_9, data_out=>output_MAC_25_9);
	MAC_25_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_10, data_out=>output_MAC_25_10);
	MAC_25_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_11, data_out=>output_MAC_25_11);
	MAC_25_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_12, data_out=>output_MAC_25_12);
	MAC_25_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_13, data_out=>output_MAC_25_13);
	MAC_25_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_14, data_out=>output_MAC_25_14);
	MAC_25_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_15, data_out=>output_MAC_25_15);
	MAC_26_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_0, data_out=>output_MAC_26_0);
	MAC_26_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_1, data_out=>output_MAC_26_1);
	MAC_26_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_2, data_out=>output_MAC_26_2);
	MAC_26_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_3, data_out=>output_MAC_26_3);
	MAC_26_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_4, data_out=>output_MAC_26_4);
	MAC_26_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_5, data_out=>output_MAC_26_5);
	MAC_26_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_6, data_out=>output_MAC_26_6);
	MAC_26_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_7, data_out=>output_MAC_26_7);
	MAC_26_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_8, data_out=>output_MAC_26_8);
	MAC_26_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_9, data_out=>output_MAC_26_9);
	MAC_26_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_10, data_out=>output_MAC_26_10);
	MAC_26_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_11, data_out=>output_MAC_26_11);
	MAC_26_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_12, data_out=>output_MAC_26_12);
	MAC_26_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_13, data_out=>output_MAC_26_13);
	MAC_26_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_14, data_out=>output_MAC_26_14);
	MAC_26_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_15, data_out=>output_MAC_26_15);
	MAC_27_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_0, data_out=>output_MAC_27_0);
	MAC_27_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_1, data_out=>output_MAC_27_1);
	MAC_27_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_2, data_out=>output_MAC_27_2);
	MAC_27_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_3, data_out=>output_MAC_27_3);
	MAC_27_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_4, data_out=>output_MAC_27_4);
	MAC_27_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_5, data_out=>output_MAC_27_5);
	MAC_27_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_6, data_out=>output_MAC_27_6);
	MAC_27_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_7, data_out=>output_MAC_27_7);
	MAC_27_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_8, data_out=>output_MAC_27_8);
	MAC_27_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_9, data_out=>output_MAC_27_9);
	MAC_27_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_10, data_out=>output_MAC_27_10);
	MAC_27_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_11, data_out=>output_MAC_27_11);
	MAC_27_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_12, data_out=>output_MAC_27_12);
	MAC_27_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_13, data_out=>output_MAC_27_13);
	MAC_27_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_14, data_out=>output_MAC_27_14);
	MAC_27_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_15, data_out=>output_MAC_27_15);
	MAC_28_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_0, data_out=>output_MAC_28_0);
	MAC_28_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_1, data_out=>output_MAC_28_1);
	MAC_28_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_2, data_out=>output_MAC_28_2);
	MAC_28_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_3, data_out=>output_MAC_28_3);
	MAC_28_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_4, data_out=>output_MAC_28_4);
	MAC_28_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_5, data_out=>output_MAC_28_5);
	MAC_28_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_6, data_out=>output_MAC_28_6);
	MAC_28_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_7, data_out=>output_MAC_28_7);
	MAC_28_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_8, data_out=>output_MAC_28_8);
	MAC_28_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_9, data_out=>output_MAC_28_9);
	MAC_28_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_10, data_out=>output_MAC_28_10);
	MAC_28_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_11, data_out=>output_MAC_28_11);
	MAC_28_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_12, data_out=>output_MAC_28_12);
	MAC_28_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_13, data_out=>output_MAC_28_13);
	MAC_28_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_14, data_out=>output_MAC_28_14);
	MAC_28_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_15, data_out=>output_MAC_28_15);
	MAC_29_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_0, data_out=>output_MAC_29_0);
	MAC_29_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_1, data_out=>output_MAC_29_1);
	MAC_29_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_2, data_out=>output_MAC_29_2);
	MAC_29_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_3, data_out=>output_MAC_29_3);
	MAC_29_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_4, data_out=>output_MAC_29_4);
	MAC_29_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_5, data_out=>output_MAC_29_5);
	MAC_29_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_6, data_out=>output_MAC_29_6);
	MAC_29_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_7, data_out=>output_MAC_29_7);
	MAC_29_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_8, data_out=>output_MAC_29_8);
	MAC_29_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_9, data_out=>output_MAC_29_9);
	MAC_29_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_10, data_out=>output_MAC_29_10);
	MAC_29_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_11, data_out=>output_MAC_29_11);
	MAC_29_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_12, data_out=>output_MAC_29_12);
	MAC_29_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_13, data_out=>output_MAC_29_13);
	MAC_29_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_14, data_out=>output_MAC_29_14);
	MAC_29_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_15, data_out=>output_MAC_29_15);
	MAC_30_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_0, data_out=>output_MAC_30_0);
	MAC_30_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_1, data_out=>output_MAC_30_1);
	MAC_30_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_2, data_out=>output_MAC_30_2);
	MAC_30_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_3, data_out=>output_MAC_30_3);
	MAC_30_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_4, data_out=>output_MAC_30_4);
	MAC_30_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_5, data_out=>output_MAC_30_5);
	MAC_30_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_6, data_out=>output_MAC_30_6);
	MAC_30_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_7, data_out=>output_MAC_30_7);
	MAC_30_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_8, data_out=>output_MAC_30_8);
	MAC_30_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_9, data_out=>output_MAC_30_9);
	MAC_30_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_10, data_out=>output_MAC_30_10);
	MAC_30_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_11, data_out=>output_MAC_30_11);
	MAC_30_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_12, data_out=>output_MAC_30_12);
	MAC_30_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_13, data_out=>output_MAC_30_13);
	MAC_30_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_14, data_out=>output_MAC_30_14);
	MAC_30_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_15, data_out=>output_MAC_30_15);
	MAC_31_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_0, data_out=>output_MAC_31_0);
	MAC_31_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_1, data_out=>output_MAC_31_1);
	MAC_31_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_2, data_out=>output_MAC_31_2);
	MAC_31_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_3, data_out=>output_MAC_31_3);
	MAC_31_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_4, data_out=>output_MAC_31_4);
	MAC_31_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_5, data_out=>output_MAC_31_5);
	MAC_31_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_6, data_out=>output_MAC_31_6);
	MAC_31_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_7, data_out=>output_MAC_31_7);
	MAC_31_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_8, data_out=>output_MAC_31_8);
	MAC_31_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_9, data_out=>output_MAC_31_9);
	MAC_31_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_10, data_out=>output_MAC_31_10);
	MAC_31_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_11, data_out=>output_MAC_31_11);
	MAC_31_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_12, data_out=>output_MAC_31_12);
	MAC_31_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_13, data_out=>output_MAC_31_13);
	MAC_31_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_14, data_out=>output_MAC_31_14);
	MAC_31_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_15, data_out=>output_MAC_31_15);

	mux_row_0: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_0_0, I1=>output_MAC_0_1, I2=>output_MAC_0_2, I3=>output_MAC_0_3, I4=>output_MAC_0_4, I5=>output_MAC_0_5, I6=>output_MAC_0_6, I7=>output_MAC_0_7, I8=>output_MAC_0_8, I9=>output_MAC_0_9, I10=>output_MAC_0_10, I11=>output_MAC_0_11, I12=>output_MAC_0_12, I13=>output_MAC_0_13, I14=>output_MAC_0_14, I15=>output_MAC_0_15, 
		SEL_mux=>SEL_mux, O=>output_row_0);

	mux_row_1: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_1_0, I1=>output_MAC_1_1, I2=>output_MAC_1_2, I3=>output_MAC_1_3, I4=>output_MAC_1_4, I5=>output_MAC_1_5, I6=>output_MAC_1_6, I7=>output_MAC_1_7, I8=>output_MAC_1_8, I9=>output_MAC_1_9, I10=>output_MAC_1_10, I11=>output_MAC_1_11, I12=>output_MAC_1_12, I13=>output_MAC_1_13, I14=>output_MAC_1_14, I15=>output_MAC_1_15, 
		SEL_mux=>SEL_mux, O=>output_row_1);

	mux_row_2: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_2_0, I1=>output_MAC_2_1, I2=>output_MAC_2_2, I3=>output_MAC_2_3, I4=>output_MAC_2_4, I5=>output_MAC_2_5, I6=>output_MAC_2_6, I7=>output_MAC_2_7, I8=>output_MAC_2_8, I9=>output_MAC_2_9, I10=>output_MAC_2_10, I11=>output_MAC_2_11, I12=>output_MAC_2_12, I13=>output_MAC_2_13, I14=>output_MAC_2_14, I15=>output_MAC_2_15, 
		SEL_mux=>SEL_mux, O=>output_row_2);

	mux_row_3: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_3_0, I1=>output_MAC_3_1, I2=>output_MAC_3_2, I3=>output_MAC_3_3, I4=>output_MAC_3_4, I5=>output_MAC_3_5, I6=>output_MAC_3_6, I7=>output_MAC_3_7, I8=>output_MAC_3_8, I9=>output_MAC_3_9, I10=>output_MAC_3_10, I11=>output_MAC_3_11, I12=>output_MAC_3_12, I13=>output_MAC_3_13, I14=>output_MAC_3_14, I15=>output_MAC_3_15, 
		SEL_mux=>SEL_mux, O=>output_row_3);

	mux_row_4: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_4_0, I1=>output_MAC_4_1, I2=>output_MAC_4_2, I3=>output_MAC_4_3, I4=>output_MAC_4_4, I5=>output_MAC_4_5, I6=>output_MAC_4_6, I7=>output_MAC_4_7, I8=>output_MAC_4_8, I9=>output_MAC_4_9, I10=>output_MAC_4_10, I11=>output_MAC_4_11, I12=>output_MAC_4_12, I13=>output_MAC_4_13, I14=>output_MAC_4_14, I15=>output_MAC_4_15, 
		SEL_mux=>SEL_mux, O=>output_row_4);

	mux_row_5: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_5_0, I1=>output_MAC_5_1, I2=>output_MAC_5_2, I3=>output_MAC_5_3, I4=>output_MAC_5_4, I5=>output_MAC_5_5, I6=>output_MAC_5_6, I7=>output_MAC_5_7, I8=>output_MAC_5_8, I9=>output_MAC_5_9, I10=>output_MAC_5_10, I11=>output_MAC_5_11, I12=>output_MAC_5_12, I13=>output_MAC_5_13, I14=>output_MAC_5_14, I15=>output_MAC_5_15, 
		SEL_mux=>SEL_mux, O=>output_row_5);

	mux_row_6: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_6_0, I1=>output_MAC_6_1, I2=>output_MAC_6_2, I3=>output_MAC_6_3, I4=>output_MAC_6_4, I5=>output_MAC_6_5, I6=>output_MAC_6_6, I7=>output_MAC_6_7, I8=>output_MAC_6_8, I9=>output_MAC_6_9, I10=>output_MAC_6_10, I11=>output_MAC_6_11, I12=>output_MAC_6_12, I13=>output_MAC_6_13, I14=>output_MAC_6_14, I15=>output_MAC_6_15, 
		SEL_mux=>SEL_mux, O=>output_row_6);

	mux_row_7: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_7_0, I1=>output_MAC_7_1, I2=>output_MAC_7_2, I3=>output_MAC_7_3, I4=>output_MAC_7_4, I5=>output_MAC_7_5, I6=>output_MAC_7_6, I7=>output_MAC_7_7, I8=>output_MAC_7_8, I9=>output_MAC_7_9, I10=>output_MAC_7_10, I11=>output_MAC_7_11, I12=>output_MAC_7_12, I13=>output_MAC_7_13, I14=>output_MAC_7_14, I15=>output_MAC_7_15, 
		SEL_mux=>SEL_mux, O=>output_row_7);

	mux_row_8: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_8_0, I1=>output_MAC_8_1, I2=>output_MAC_8_2, I3=>output_MAC_8_3, I4=>output_MAC_8_4, I5=>output_MAC_8_5, I6=>output_MAC_8_6, I7=>output_MAC_8_7, I8=>output_MAC_8_8, I9=>output_MAC_8_9, I10=>output_MAC_8_10, I11=>output_MAC_8_11, I12=>output_MAC_8_12, I13=>output_MAC_8_13, I14=>output_MAC_8_14, I15=>output_MAC_8_15, 
		SEL_mux=>SEL_mux, O=>output_row_8);

	mux_row_9: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_9_0, I1=>output_MAC_9_1, I2=>output_MAC_9_2, I3=>output_MAC_9_3, I4=>output_MAC_9_4, I5=>output_MAC_9_5, I6=>output_MAC_9_6, I7=>output_MAC_9_7, I8=>output_MAC_9_8, I9=>output_MAC_9_9, I10=>output_MAC_9_10, I11=>output_MAC_9_11, I12=>output_MAC_9_12, I13=>output_MAC_9_13, I14=>output_MAC_9_14, I15=>output_MAC_9_15, 
		SEL_mux=>SEL_mux, O=>output_row_9);

	mux_row_10: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_10_0, I1=>output_MAC_10_1, I2=>output_MAC_10_2, I3=>output_MAC_10_3, I4=>output_MAC_10_4, I5=>output_MAC_10_5, I6=>output_MAC_10_6, I7=>output_MAC_10_7, I8=>output_MAC_10_8, I9=>output_MAC_10_9, I10=>output_MAC_10_10, I11=>output_MAC_10_11, I12=>output_MAC_10_12, I13=>output_MAC_10_13, I14=>output_MAC_10_14, I15=>output_MAC_10_15, 
		SEL_mux=>SEL_mux, O=>output_row_10);

	mux_row_11: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_11_0, I1=>output_MAC_11_1, I2=>output_MAC_11_2, I3=>output_MAC_11_3, I4=>output_MAC_11_4, I5=>output_MAC_11_5, I6=>output_MAC_11_6, I7=>output_MAC_11_7, I8=>output_MAC_11_8, I9=>output_MAC_11_9, I10=>output_MAC_11_10, I11=>output_MAC_11_11, I12=>output_MAC_11_12, I13=>output_MAC_11_13, I14=>output_MAC_11_14, I15=>output_MAC_11_15, 
		SEL_mux=>SEL_mux, O=>output_row_11);

	mux_row_12: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_12_0, I1=>output_MAC_12_1, I2=>output_MAC_12_2, I3=>output_MAC_12_3, I4=>output_MAC_12_4, I5=>output_MAC_12_5, I6=>output_MAC_12_6, I7=>output_MAC_12_7, I8=>output_MAC_12_8, I9=>output_MAC_12_9, I10=>output_MAC_12_10, I11=>output_MAC_12_11, I12=>output_MAC_12_12, I13=>output_MAC_12_13, I14=>output_MAC_12_14, I15=>output_MAC_12_15, 
		SEL_mux=>SEL_mux, O=>output_row_12);

	mux_row_13: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_13_0, I1=>output_MAC_13_1, I2=>output_MAC_13_2, I3=>output_MAC_13_3, I4=>output_MAC_13_4, I5=>output_MAC_13_5, I6=>output_MAC_13_6, I7=>output_MAC_13_7, I8=>output_MAC_13_8, I9=>output_MAC_13_9, I10=>output_MAC_13_10, I11=>output_MAC_13_11, I12=>output_MAC_13_12, I13=>output_MAC_13_13, I14=>output_MAC_13_14, I15=>output_MAC_13_15, 
		SEL_mux=>SEL_mux, O=>output_row_13);

	mux_row_14: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_14_0, I1=>output_MAC_14_1, I2=>output_MAC_14_2, I3=>output_MAC_14_3, I4=>output_MAC_14_4, I5=>output_MAC_14_5, I6=>output_MAC_14_6, I7=>output_MAC_14_7, I8=>output_MAC_14_8, I9=>output_MAC_14_9, I10=>output_MAC_14_10, I11=>output_MAC_14_11, I12=>output_MAC_14_12, I13=>output_MAC_14_13, I14=>output_MAC_14_14, I15=>output_MAC_14_15, 
		SEL_mux=>SEL_mux, O=>output_row_14);

	mux_row_15: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_15_0, I1=>output_MAC_15_1, I2=>output_MAC_15_2, I3=>output_MAC_15_3, I4=>output_MAC_15_4, I5=>output_MAC_15_5, I6=>output_MAC_15_6, I7=>output_MAC_15_7, I8=>output_MAC_15_8, I9=>output_MAC_15_9, I10=>output_MAC_15_10, I11=>output_MAC_15_11, I12=>output_MAC_15_12, I13=>output_MAC_15_13, I14=>output_MAC_15_14, I15=>output_MAC_15_15, 
		SEL_mux=>SEL_mux, O=>output_row_15);

	mux_row_16: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_16_0, I1=>output_MAC_16_1, I2=>output_MAC_16_2, I3=>output_MAC_16_3, I4=>output_MAC_16_4, I5=>output_MAC_16_5, I6=>output_MAC_16_6, I7=>output_MAC_16_7, I8=>output_MAC_16_8, I9=>output_MAC_16_9, I10=>output_MAC_16_10, I11=>output_MAC_16_11, I12=>output_MAC_16_12, I13=>output_MAC_16_13, I14=>output_MAC_16_14, I15=>output_MAC_16_15, 
		SEL_mux=>SEL_mux, O=>output_row_16);

	mux_row_17: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_17_0, I1=>output_MAC_17_1, I2=>output_MAC_17_2, I3=>output_MAC_17_3, I4=>output_MAC_17_4, I5=>output_MAC_17_5, I6=>output_MAC_17_6, I7=>output_MAC_17_7, I8=>output_MAC_17_8, I9=>output_MAC_17_9, I10=>output_MAC_17_10, I11=>output_MAC_17_11, I12=>output_MAC_17_12, I13=>output_MAC_17_13, I14=>output_MAC_17_14, I15=>output_MAC_17_15, 
		SEL_mux=>SEL_mux, O=>output_row_17);

	mux_row_18: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_18_0, I1=>output_MAC_18_1, I2=>output_MAC_18_2, I3=>output_MAC_18_3, I4=>output_MAC_18_4, I5=>output_MAC_18_5, I6=>output_MAC_18_6, I7=>output_MAC_18_7, I8=>output_MAC_18_8, I9=>output_MAC_18_9, I10=>output_MAC_18_10, I11=>output_MAC_18_11, I12=>output_MAC_18_12, I13=>output_MAC_18_13, I14=>output_MAC_18_14, I15=>output_MAC_18_15, 
		SEL_mux=>SEL_mux, O=>output_row_18);

	mux_row_19: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_19_0, I1=>output_MAC_19_1, I2=>output_MAC_19_2, I3=>output_MAC_19_3, I4=>output_MAC_19_4, I5=>output_MAC_19_5, I6=>output_MAC_19_6, I7=>output_MAC_19_7, I8=>output_MAC_19_8, I9=>output_MAC_19_9, I10=>output_MAC_19_10, I11=>output_MAC_19_11, I12=>output_MAC_19_12, I13=>output_MAC_19_13, I14=>output_MAC_19_14, I15=>output_MAC_19_15, 
		SEL_mux=>SEL_mux, O=>output_row_19);

	mux_row_20: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_20_0, I1=>output_MAC_20_1, I2=>output_MAC_20_2, I3=>output_MAC_20_3, I4=>output_MAC_20_4, I5=>output_MAC_20_5, I6=>output_MAC_20_6, I7=>output_MAC_20_7, I8=>output_MAC_20_8, I9=>output_MAC_20_9, I10=>output_MAC_20_10, I11=>output_MAC_20_11, I12=>output_MAC_20_12, I13=>output_MAC_20_13, I14=>output_MAC_20_14, I15=>output_MAC_20_15, 
		SEL_mux=>SEL_mux, O=>output_row_20);

	mux_row_21: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_21_0, I1=>output_MAC_21_1, I2=>output_MAC_21_2, I3=>output_MAC_21_3, I4=>output_MAC_21_4, I5=>output_MAC_21_5, I6=>output_MAC_21_6, I7=>output_MAC_21_7, I8=>output_MAC_21_8, I9=>output_MAC_21_9, I10=>output_MAC_21_10, I11=>output_MAC_21_11, I12=>output_MAC_21_12, I13=>output_MAC_21_13, I14=>output_MAC_21_14, I15=>output_MAC_21_15, 
		SEL_mux=>SEL_mux, O=>output_row_21);

	mux_row_22: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_22_0, I1=>output_MAC_22_1, I2=>output_MAC_22_2, I3=>output_MAC_22_3, I4=>output_MAC_22_4, I5=>output_MAC_22_5, I6=>output_MAC_22_6, I7=>output_MAC_22_7, I8=>output_MAC_22_8, I9=>output_MAC_22_9, I10=>output_MAC_22_10, I11=>output_MAC_22_11, I12=>output_MAC_22_12, I13=>output_MAC_22_13, I14=>output_MAC_22_14, I15=>output_MAC_22_15, 
		SEL_mux=>SEL_mux, O=>output_row_22);

	mux_row_23: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_23_0, I1=>output_MAC_23_1, I2=>output_MAC_23_2, I3=>output_MAC_23_3, I4=>output_MAC_23_4, I5=>output_MAC_23_5, I6=>output_MAC_23_6, I7=>output_MAC_23_7, I8=>output_MAC_23_8, I9=>output_MAC_23_9, I10=>output_MAC_23_10, I11=>output_MAC_23_11, I12=>output_MAC_23_12, I13=>output_MAC_23_13, I14=>output_MAC_23_14, I15=>output_MAC_23_15, 
		SEL_mux=>SEL_mux, O=>output_row_23);

	mux_row_24: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_24_0, I1=>output_MAC_24_1, I2=>output_MAC_24_2, I3=>output_MAC_24_3, I4=>output_MAC_24_4, I5=>output_MAC_24_5, I6=>output_MAC_24_6, I7=>output_MAC_24_7, I8=>output_MAC_24_8, I9=>output_MAC_24_9, I10=>output_MAC_24_10, I11=>output_MAC_24_11, I12=>output_MAC_24_12, I13=>output_MAC_24_13, I14=>output_MAC_24_14, I15=>output_MAC_24_15, 
		SEL_mux=>SEL_mux, O=>output_row_24);

	mux_row_25: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_25_0, I1=>output_MAC_25_1, I2=>output_MAC_25_2, I3=>output_MAC_25_3, I4=>output_MAC_25_4, I5=>output_MAC_25_5, I6=>output_MAC_25_6, I7=>output_MAC_25_7, I8=>output_MAC_25_8, I9=>output_MAC_25_9, I10=>output_MAC_25_10, I11=>output_MAC_25_11, I12=>output_MAC_25_12, I13=>output_MAC_25_13, I14=>output_MAC_25_14, I15=>output_MAC_25_15, 
		SEL_mux=>SEL_mux, O=>output_row_25);

	mux_row_26: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_26_0, I1=>output_MAC_26_1, I2=>output_MAC_26_2, I3=>output_MAC_26_3, I4=>output_MAC_26_4, I5=>output_MAC_26_5, I6=>output_MAC_26_6, I7=>output_MAC_26_7, I8=>output_MAC_26_8, I9=>output_MAC_26_9, I10=>output_MAC_26_10, I11=>output_MAC_26_11, I12=>output_MAC_26_12, I13=>output_MAC_26_13, I14=>output_MAC_26_14, I15=>output_MAC_26_15, 
		SEL_mux=>SEL_mux, O=>output_row_26);

	mux_row_27: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_27_0, I1=>output_MAC_27_1, I2=>output_MAC_27_2, I3=>output_MAC_27_3, I4=>output_MAC_27_4, I5=>output_MAC_27_5, I6=>output_MAC_27_6, I7=>output_MAC_27_7, I8=>output_MAC_27_8, I9=>output_MAC_27_9, I10=>output_MAC_27_10, I11=>output_MAC_27_11, I12=>output_MAC_27_12, I13=>output_MAC_27_13, I14=>output_MAC_27_14, I15=>output_MAC_27_15, 
		SEL_mux=>SEL_mux, O=>output_row_27);

	mux_row_28: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_28_0, I1=>output_MAC_28_1, I2=>output_MAC_28_2, I3=>output_MAC_28_3, I4=>output_MAC_28_4, I5=>output_MAC_28_5, I6=>output_MAC_28_6, I7=>output_MAC_28_7, I8=>output_MAC_28_8, I9=>output_MAC_28_9, I10=>output_MAC_28_10, I11=>output_MAC_28_11, I12=>output_MAC_28_12, I13=>output_MAC_28_13, I14=>output_MAC_28_14, I15=>output_MAC_28_15, 
		SEL_mux=>SEL_mux, O=>output_row_28);

	mux_row_29: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_29_0, I1=>output_MAC_29_1, I2=>output_MAC_29_2, I3=>output_MAC_29_3, I4=>output_MAC_29_4, I5=>output_MAC_29_5, I6=>output_MAC_29_6, I7=>output_MAC_29_7, I8=>output_MAC_29_8, I9=>output_MAC_29_9, I10=>output_MAC_29_10, I11=>output_MAC_29_11, I12=>output_MAC_29_12, I13=>output_MAC_29_13, I14=>output_MAC_29_14, I15=>output_MAC_29_15, 
		SEL_mux=>SEL_mux, O=>output_row_29);

	mux_row_30: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_30_0, I1=>output_MAC_30_1, I2=>output_MAC_30_2, I3=>output_MAC_30_3, I4=>output_MAC_30_4, I5=>output_MAC_30_5, I6=>output_MAC_30_6, I7=>output_MAC_30_7, I8=>output_MAC_30_8, I9=>output_MAC_30_9, I10=>output_MAC_30_10, I11=>output_MAC_30_11, I12=>output_MAC_30_12, I13=>output_MAC_30_13, I14=>output_MAC_30_14, I15=>output_MAC_30_15, 
		SEL_mux=>SEL_mux, O=>output_row_30);

	mux_row_31: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_31_0, I1=>output_MAC_31_1, I2=>output_MAC_31_2, I3=>output_MAC_31_3, I4=>output_MAC_31_4, I5=>output_MAC_31_5, I6=>output_MAC_31_6, I7=>output_MAC_31_7, I8=>output_MAC_31_8, I9=>output_MAC_31_9, I10=>output_MAC_31_10, I11=>output_MAC_31_11, I12=>output_MAC_31_12, I13=>output_MAC_31_13, I14=>output_MAC_31_14, I15=>output_MAC_31_15, 
		SEL_mux=>SEL_mux, O=>output_row_31);


END behaviour;
