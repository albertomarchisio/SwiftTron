
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MAC_64x32_8 IS
PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7, input_row_8, input_row_9, 
	input_row_10, input_row_11, input_row_12, input_row_13, input_row_14, input_row_15, input_row_16, input_row_17, input_row_18, input_row_19, 
	input_row_20, input_row_21, input_row_22, input_row_23, input_row_24, input_row_25, input_row_26, input_row_27, input_row_28, input_row_29, 
	input_row_30, input_row_31, input_row_32, input_row_33, input_row_34, input_row_35, input_row_36, input_row_37, input_row_38, input_row_39, 
	input_row_40, input_row_41, input_row_42, input_row_43, input_row_44, input_row_45, input_row_46, input_row_47, input_row_48, input_row_49, 
	input_row_50, input_row_51, input_row_52, input_row_53, input_row_54, input_row_55, input_row_56, input_row_57, input_row_58, input_row_59, 
	input_row_60, input_row_61, input_row_62, input_row_63: IN STD_LOGIC_VECTOR(7 downto 0);
	input_col_0, input_col_1, input_col_2, input_col_3, input_col_4, input_col_5, input_col_6, input_col_7, input_col_8, input_col_9, 
	input_col_10, input_col_11, input_col_12, input_col_13, input_col_14, input_col_15, input_col_16, input_col_17, input_col_18, input_col_19, 
	input_col_20, input_col_21, input_col_22, input_col_23, input_col_24, input_col_25, input_col_26, input_col_27, input_col_28, input_col_29, 
	input_col_30, input_col_31: IN STD_LOGIC_VECTOR(7 downto 0);
	SEL_mux: IN STD_LOGIC_VECTOR(4 downto 0);
	CLK, RST_n, ENABLE : IN STD_LOGIC;
	output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7, output_row_8, output_row_9, 
	output_row_10, output_row_11, output_row_12, output_row_13, output_row_14, output_row_15, output_row_16, output_row_17, output_row_18, output_row_19, 
	output_row_20, output_row_21, output_row_22, output_row_23, output_row_24, output_row_25, output_row_26, output_row_27, output_row_28, output_row_29, 
	output_row_30, output_row_31, output_row_32, output_row_33, output_row_34, output_row_35, output_row_36, output_row_37, output_row_38, output_row_39, 
	output_row_40, output_row_41, output_row_42, output_row_43, output_row_44, output_row_45, output_row_46, output_row_47, output_row_48, output_row_49, 
	output_row_50, output_row_51, output_row_52, output_row_53, output_row_54, output_row_55, output_row_56, output_row_57, output_row_58, output_row_59, 
	output_row_60, output_row_61, output_row_62, output_row_63: OUT STD_LOGIC_VECTOR(31 downto 0)
);
END MAC_64x32_8;

ARCHITECTURE behaviour OF  MAC_64x32_8 IS

	COMPONENT MAC IS
	GENERIC (data_size : POSITIVE := 2;
	 acc_size : POSITIVE := 16 );
	PORT( data_in_A, data_in_B  : IN STD_LOGIC_VECTOR(data_size-1 downto 0);
		CLK, RST_n, ENABLE 	: IN STD_LOGIC;
		data_out    			: OUT STD_LOGIC_VECTOR(acc_size-1 downto 0));
	END COMPONENT;

	COMPONENT mux_32to1_nbit IS
	GENERIC ( N : POSITIVE :=2);
	PORT(
		I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, 
		I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, 
		I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, 
		I30, I31: IN STD_LOGIC_VECTOR(N-1 downto 0);
		SEL_mux  : IN STD_LOGIC_VECTOR(4 downto 0);
		O    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
	END COMPONENT;


	SIGNAL output_MAC_0_0, output_MAC_0_1, output_MAC_0_2, output_MAC_0_3, output_MAC_0_4, output_MAC_0_5, output_MAC_0_6, output_MAC_0_7, output_MAC_0_8, output_MAC_0_9, 
		output_MAC_0_10, output_MAC_0_11, output_MAC_0_12, output_MAC_0_13, output_MAC_0_14, output_MAC_0_15, output_MAC_0_16, output_MAC_0_17, output_MAC_0_18, output_MAC_0_19, 
		output_MAC_0_20, output_MAC_0_21, output_MAC_0_22, output_MAC_0_23, output_MAC_0_24, output_MAC_0_25, output_MAC_0_26, output_MAC_0_27, output_MAC_0_28, output_MAC_0_29, 
		output_MAC_0_30, output_MAC_0_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_1_0, output_MAC_1_1, output_MAC_1_2, output_MAC_1_3, output_MAC_1_4, output_MAC_1_5, output_MAC_1_6, output_MAC_1_7, output_MAC_1_8, output_MAC_1_9, 
		output_MAC_1_10, output_MAC_1_11, output_MAC_1_12, output_MAC_1_13, output_MAC_1_14, output_MAC_1_15, output_MAC_1_16, output_MAC_1_17, output_MAC_1_18, output_MAC_1_19, 
		output_MAC_1_20, output_MAC_1_21, output_MAC_1_22, output_MAC_1_23, output_MAC_1_24, output_MAC_1_25, output_MAC_1_26, output_MAC_1_27, output_MAC_1_28, output_MAC_1_29, 
		output_MAC_1_30, output_MAC_1_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_2_0, output_MAC_2_1, output_MAC_2_2, output_MAC_2_3, output_MAC_2_4, output_MAC_2_5, output_MAC_2_6, output_MAC_2_7, output_MAC_2_8, output_MAC_2_9, 
		output_MAC_2_10, output_MAC_2_11, output_MAC_2_12, output_MAC_2_13, output_MAC_2_14, output_MAC_2_15, output_MAC_2_16, output_MAC_2_17, output_MAC_2_18, output_MAC_2_19, 
		output_MAC_2_20, output_MAC_2_21, output_MAC_2_22, output_MAC_2_23, output_MAC_2_24, output_MAC_2_25, output_MAC_2_26, output_MAC_2_27, output_MAC_2_28, output_MAC_2_29, 
		output_MAC_2_30, output_MAC_2_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_3_0, output_MAC_3_1, output_MAC_3_2, output_MAC_3_3, output_MAC_3_4, output_MAC_3_5, output_MAC_3_6, output_MAC_3_7, output_MAC_3_8, output_MAC_3_9, 
		output_MAC_3_10, output_MAC_3_11, output_MAC_3_12, output_MAC_3_13, output_MAC_3_14, output_MAC_3_15, output_MAC_3_16, output_MAC_3_17, output_MAC_3_18, output_MAC_3_19, 
		output_MAC_3_20, output_MAC_3_21, output_MAC_3_22, output_MAC_3_23, output_MAC_3_24, output_MAC_3_25, output_MAC_3_26, output_MAC_3_27, output_MAC_3_28, output_MAC_3_29, 
		output_MAC_3_30, output_MAC_3_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_4_0, output_MAC_4_1, output_MAC_4_2, output_MAC_4_3, output_MAC_4_4, output_MAC_4_5, output_MAC_4_6, output_MAC_4_7, output_MAC_4_8, output_MAC_4_9, 
		output_MAC_4_10, output_MAC_4_11, output_MAC_4_12, output_MAC_4_13, output_MAC_4_14, output_MAC_4_15, output_MAC_4_16, output_MAC_4_17, output_MAC_4_18, output_MAC_4_19, 
		output_MAC_4_20, output_MAC_4_21, output_MAC_4_22, output_MAC_4_23, output_MAC_4_24, output_MAC_4_25, output_MAC_4_26, output_MAC_4_27, output_MAC_4_28, output_MAC_4_29, 
		output_MAC_4_30, output_MAC_4_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_5_0, output_MAC_5_1, output_MAC_5_2, output_MAC_5_3, output_MAC_5_4, output_MAC_5_5, output_MAC_5_6, output_MAC_5_7, output_MAC_5_8, output_MAC_5_9, 
		output_MAC_5_10, output_MAC_5_11, output_MAC_5_12, output_MAC_5_13, output_MAC_5_14, output_MAC_5_15, output_MAC_5_16, output_MAC_5_17, output_MAC_5_18, output_MAC_5_19, 
		output_MAC_5_20, output_MAC_5_21, output_MAC_5_22, output_MAC_5_23, output_MAC_5_24, output_MAC_5_25, output_MAC_5_26, output_MAC_5_27, output_MAC_5_28, output_MAC_5_29, 
		output_MAC_5_30, output_MAC_5_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_6_0, output_MAC_6_1, output_MAC_6_2, output_MAC_6_3, output_MAC_6_4, output_MAC_6_5, output_MAC_6_6, output_MAC_6_7, output_MAC_6_8, output_MAC_6_9, 
		output_MAC_6_10, output_MAC_6_11, output_MAC_6_12, output_MAC_6_13, output_MAC_6_14, output_MAC_6_15, output_MAC_6_16, output_MAC_6_17, output_MAC_6_18, output_MAC_6_19, 
		output_MAC_6_20, output_MAC_6_21, output_MAC_6_22, output_MAC_6_23, output_MAC_6_24, output_MAC_6_25, output_MAC_6_26, output_MAC_6_27, output_MAC_6_28, output_MAC_6_29, 
		output_MAC_6_30, output_MAC_6_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_7_0, output_MAC_7_1, output_MAC_7_2, output_MAC_7_3, output_MAC_7_4, output_MAC_7_5, output_MAC_7_6, output_MAC_7_7, output_MAC_7_8, output_MAC_7_9, 
		output_MAC_7_10, output_MAC_7_11, output_MAC_7_12, output_MAC_7_13, output_MAC_7_14, output_MAC_7_15, output_MAC_7_16, output_MAC_7_17, output_MAC_7_18, output_MAC_7_19, 
		output_MAC_7_20, output_MAC_7_21, output_MAC_7_22, output_MAC_7_23, output_MAC_7_24, output_MAC_7_25, output_MAC_7_26, output_MAC_7_27, output_MAC_7_28, output_MAC_7_29, 
		output_MAC_7_30, output_MAC_7_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_8_0, output_MAC_8_1, output_MAC_8_2, output_MAC_8_3, output_MAC_8_4, output_MAC_8_5, output_MAC_8_6, output_MAC_8_7, output_MAC_8_8, output_MAC_8_9, 
		output_MAC_8_10, output_MAC_8_11, output_MAC_8_12, output_MAC_8_13, output_MAC_8_14, output_MAC_8_15, output_MAC_8_16, output_MAC_8_17, output_MAC_8_18, output_MAC_8_19, 
		output_MAC_8_20, output_MAC_8_21, output_MAC_8_22, output_MAC_8_23, output_MAC_8_24, output_MAC_8_25, output_MAC_8_26, output_MAC_8_27, output_MAC_8_28, output_MAC_8_29, 
		output_MAC_8_30, output_MAC_8_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_9_0, output_MAC_9_1, output_MAC_9_2, output_MAC_9_3, output_MAC_9_4, output_MAC_9_5, output_MAC_9_6, output_MAC_9_7, output_MAC_9_8, output_MAC_9_9, 
		output_MAC_9_10, output_MAC_9_11, output_MAC_9_12, output_MAC_9_13, output_MAC_9_14, output_MAC_9_15, output_MAC_9_16, output_MAC_9_17, output_MAC_9_18, output_MAC_9_19, 
		output_MAC_9_20, output_MAC_9_21, output_MAC_9_22, output_MAC_9_23, output_MAC_9_24, output_MAC_9_25, output_MAC_9_26, output_MAC_9_27, output_MAC_9_28, output_MAC_9_29, 
		output_MAC_9_30, output_MAC_9_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_10_0, output_MAC_10_1, output_MAC_10_2, output_MAC_10_3, output_MAC_10_4, output_MAC_10_5, output_MAC_10_6, output_MAC_10_7, output_MAC_10_8, output_MAC_10_9, 
		output_MAC_10_10, output_MAC_10_11, output_MAC_10_12, output_MAC_10_13, output_MAC_10_14, output_MAC_10_15, output_MAC_10_16, output_MAC_10_17, output_MAC_10_18, output_MAC_10_19, 
		output_MAC_10_20, output_MAC_10_21, output_MAC_10_22, output_MAC_10_23, output_MAC_10_24, output_MAC_10_25, output_MAC_10_26, output_MAC_10_27, output_MAC_10_28, output_MAC_10_29, 
		output_MAC_10_30, output_MAC_10_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_11_0, output_MAC_11_1, output_MAC_11_2, output_MAC_11_3, output_MAC_11_4, output_MAC_11_5, output_MAC_11_6, output_MAC_11_7, output_MAC_11_8, output_MAC_11_9, 
		output_MAC_11_10, output_MAC_11_11, output_MAC_11_12, output_MAC_11_13, output_MAC_11_14, output_MAC_11_15, output_MAC_11_16, output_MAC_11_17, output_MAC_11_18, output_MAC_11_19, 
		output_MAC_11_20, output_MAC_11_21, output_MAC_11_22, output_MAC_11_23, output_MAC_11_24, output_MAC_11_25, output_MAC_11_26, output_MAC_11_27, output_MAC_11_28, output_MAC_11_29, 
		output_MAC_11_30, output_MAC_11_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_12_0, output_MAC_12_1, output_MAC_12_2, output_MAC_12_3, output_MAC_12_4, output_MAC_12_5, output_MAC_12_6, output_MAC_12_7, output_MAC_12_8, output_MAC_12_9, 
		output_MAC_12_10, output_MAC_12_11, output_MAC_12_12, output_MAC_12_13, output_MAC_12_14, output_MAC_12_15, output_MAC_12_16, output_MAC_12_17, output_MAC_12_18, output_MAC_12_19, 
		output_MAC_12_20, output_MAC_12_21, output_MAC_12_22, output_MAC_12_23, output_MAC_12_24, output_MAC_12_25, output_MAC_12_26, output_MAC_12_27, output_MAC_12_28, output_MAC_12_29, 
		output_MAC_12_30, output_MAC_12_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_13_0, output_MAC_13_1, output_MAC_13_2, output_MAC_13_3, output_MAC_13_4, output_MAC_13_5, output_MAC_13_6, output_MAC_13_7, output_MAC_13_8, output_MAC_13_9, 
		output_MAC_13_10, output_MAC_13_11, output_MAC_13_12, output_MAC_13_13, output_MAC_13_14, output_MAC_13_15, output_MAC_13_16, output_MAC_13_17, output_MAC_13_18, output_MAC_13_19, 
		output_MAC_13_20, output_MAC_13_21, output_MAC_13_22, output_MAC_13_23, output_MAC_13_24, output_MAC_13_25, output_MAC_13_26, output_MAC_13_27, output_MAC_13_28, output_MAC_13_29, 
		output_MAC_13_30, output_MAC_13_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_14_0, output_MAC_14_1, output_MAC_14_2, output_MAC_14_3, output_MAC_14_4, output_MAC_14_5, output_MAC_14_6, output_MAC_14_7, output_MAC_14_8, output_MAC_14_9, 
		output_MAC_14_10, output_MAC_14_11, output_MAC_14_12, output_MAC_14_13, output_MAC_14_14, output_MAC_14_15, output_MAC_14_16, output_MAC_14_17, output_MAC_14_18, output_MAC_14_19, 
		output_MAC_14_20, output_MAC_14_21, output_MAC_14_22, output_MAC_14_23, output_MAC_14_24, output_MAC_14_25, output_MAC_14_26, output_MAC_14_27, output_MAC_14_28, output_MAC_14_29, 
		output_MAC_14_30, output_MAC_14_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_15_0, output_MAC_15_1, output_MAC_15_2, output_MAC_15_3, output_MAC_15_4, output_MAC_15_5, output_MAC_15_6, output_MAC_15_7, output_MAC_15_8, output_MAC_15_9, 
		output_MAC_15_10, output_MAC_15_11, output_MAC_15_12, output_MAC_15_13, output_MAC_15_14, output_MAC_15_15, output_MAC_15_16, output_MAC_15_17, output_MAC_15_18, output_MAC_15_19, 
		output_MAC_15_20, output_MAC_15_21, output_MAC_15_22, output_MAC_15_23, output_MAC_15_24, output_MAC_15_25, output_MAC_15_26, output_MAC_15_27, output_MAC_15_28, output_MAC_15_29, 
		output_MAC_15_30, output_MAC_15_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_16_0, output_MAC_16_1, output_MAC_16_2, output_MAC_16_3, output_MAC_16_4, output_MAC_16_5, output_MAC_16_6, output_MAC_16_7, output_MAC_16_8, output_MAC_16_9, 
		output_MAC_16_10, output_MAC_16_11, output_MAC_16_12, output_MAC_16_13, output_MAC_16_14, output_MAC_16_15, output_MAC_16_16, output_MAC_16_17, output_MAC_16_18, output_MAC_16_19, 
		output_MAC_16_20, output_MAC_16_21, output_MAC_16_22, output_MAC_16_23, output_MAC_16_24, output_MAC_16_25, output_MAC_16_26, output_MAC_16_27, output_MAC_16_28, output_MAC_16_29, 
		output_MAC_16_30, output_MAC_16_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_17_0, output_MAC_17_1, output_MAC_17_2, output_MAC_17_3, output_MAC_17_4, output_MAC_17_5, output_MAC_17_6, output_MAC_17_7, output_MAC_17_8, output_MAC_17_9, 
		output_MAC_17_10, output_MAC_17_11, output_MAC_17_12, output_MAC_17_13, output_MAC_17_14, output_MAC_17_15, output_MAC_17_16, output_MAC_17_17, output_MAC_17_18, output_MAC_17_19, 
		output_MAC_17_20, output_MAC_17_21, output_MAC_17_22, output_MAC_17_23, output_MAC_17_24, output_MAC_17_25, output_MAC_17_26, output_MAC_17_27, output_MAC_17_28, output_MAC_17_29, 
		output_MAC_17_30, output_MAC_17_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_18_0, output_MAC_18_1, output_MAC_18_2, output_MAC_18_3, output_MAC_18_4, output_MAC_18_5, output_MAC_18_6, output_MAC_18_7, output_MAC_18_8, output_MAC_18_9, 
		output_MAC_18_10, output_MAC_18_11, output_MAC_18_12, output_MAC_18_13, output_MAC_18_14, output_MAC_18_15, output_MAC_18_16, output_MAC_18_17, output_MAC_18_18, output_MAC_18_19, 
		output_MAC_18_20, output_MAC_18_21, output_MAC_18_22, output_MAC_18_23, output_MAC_18_24, output_MAC_18_25, output_MAC_18_26, output_MAC_18_27, output_MAC_18_28, output_MAC_18_29, 
		output_MAC_18_30, output_MAC_18_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_19_0, output_MAC_19_1, output_MAC_19_2, output_MAC_19_3, output_MAC_19_4, output_MAC_19_5, output_MAC_19_6, output_MAC_19_7, output_MAC_19_8, output_MAC_19_9, 
		output_MAC_19_10, output_MAC_19_11, output_MAC_19_12, output_MAC_19_13, output_MAC_19_14, output_MAC_19_15, output_MAC_19_16, output_MAC_19_17, output_MAC_19_18, output_MAC_19_19, 
		output_MAC_19_20, output_MAC_19_21, output_MAC_19_22, output_MAC_19_23, output_MAC_19_24, output_MAC_19_25, output_MAC_19_26, output_MAC_19_27, output_MAC_19_28, output_MAC_19_29, 
		output_MAC_19_30, output_MAC_19_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_20_0, output_MAC_20_1, output_MAC_20_2, output_MAC_20_3, output_MAC_20_4, output_MAC_20_5, output_MAC_20_6, output_MAC_20_7, output_MAC_20_8, output_MAC_20_9, 
		output_MAC_20_10, output_MAC_20_11, output_MAC_20_12, output_MAC_20_13, output_MAC_20_14, output_MAC_20_15, output_MAC_20_16, output_MAC_20_17, output_MAC_20_18, output_MAC_20_19, 
		output_MAC_20_20, output_MAC_20_21, output_MAC_20_22, output_MAC_20_23, output_MAC_20_24, output_MAC_20_25, output_MAC_20_26, output_MAC_20_27, output_MAC_20_28, output_MAC_20_29, 
		output_MAC_20_30, output_MAC_20_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_21_0, output_MAC_21_1, output_MAC_21_2, output_MAC_21_3, output_MAC_21_4, output_MAC_21_5, output_MAC_21_6, output_MAC_21_7, output_MAC_21_8, output_MAC_21_9, 
		output_MAC_21_10, output_MAC_21_11, output_MAC_21_12, output_MAC_21_13, output_MAC_21_14, output_MAC_21_15, output_MAC_21_16, output_MAC_21_17, output_MAC_21_18, output_MAC_21_19, 
		output_MAC_21_20, output_MAC_21_21, output_MAC_21_22, output_MAC_21_23, output_MAC_21_24, output_MAC_21_25, output_MAC_21_26, output_MAC_21_27, output_MAC_21_28, output_MAC_21_29, 
		output_MAC_21_30, output_MAC_21_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_22_0, output_MAC_22_1, output_MAC_22_2, output_MAC_22_3, output_MAC_22_4, output_MAC_22_5, output_MAC_22_6, output_MAC_22_7, output_MAC_22_8, output_MAC_22_9, 
		output_MAC_22_10, output_MAC_22_11, output_MAC_22_12, output_MAC_22_13, output_MAC_22_14, output_MAC_22_15, output_MAC_22_16, output_MAC_22_17, output_MAC_22_18, output_MAC_22_19, 
		output_MAC_22_20, output_MAC_22_21, output_MAC_22_22, output_MAC_22_23, output_MAC_22_24, output_MAC_22_25, output_MAC_22_26, output_MAC_22_27, output_MAC_22_28, output_MAC_22_29, 
		output_MAC_22_30, output_MAC_22_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_23_0, output_MAC_23_1, output_MAC_23_2, output_MAC_23_3, output_MAC_23_4, output_MAC_23_5, output_MAC_23_6, output_MAC_23_7, output_MAC_23_8, output_MAC_23_9, 
		output_MAC_23_10, output_MAC_23_11, output_MAC_23_12, output_MAC_23_13, output_MAC_23_14, output_MAC_23_15, output_MAC_23_16, output_MAC_23_17, output_MAC_23_18, output_MAC_23_19, 
		output_MAC_23_20, output_MAC_23_21, output_MAC_23_22, output_MAC_23_23, output_MAC_23_24, output_MAC_23_25, output_MAC_23_26, output_MAC_23_27, output_MAC_23_28, output_MAC_23_29, 
		output_MAC_23_30, output_MAC_23_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_24_0, output_MAC_24_1, output_MAC_24_2, output_MAC_24_3, output_MAC_24_4, output_MAC_24_5, output_MAC_24_6, output_MAC_24_7, output_MAC_24_8, output_MAC_24_9, 
		output_MAC_24_10, output_MAC_24_11, output_MAC_24_12, output_MAC_24_13, output_MAC_24_14, output_MAC_24_15, output_MAC_24_16, output_MAC_24_17, output_MAC_24_18, output_MAC_24_19, 
		output_MAC_24_20, output_MAC_24_21, output_MAC_24_22, output_MAC_24_23, output_MAC_24_24, output_MAC_24_25, output_MAC_24_26, output_MAC_24_27, output_MAC_24_28, output_MAC_24_29, 
		output_MAC_24_30, output_MAC_24_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_25_0, output_MAC_25_1, output_MAC_25_2, output_MAC_25_3, output_MAC_25_4, output_MAC_25_5, output_MAC_25_6, output_MAC_25_7, output_MAC_25_8, output_MAC_25_9, 
		output_MAC_25_10, output_MAC_25_11, output_MAC_25_12, output_MAC_25_13, output_MAC_25_14, output_MAC_25_15, output_MAC_25_16, output_MAC_25_17, output_MAC_25_18, output_MAC_25_19, 
		output_MAC_25_20, output_MAC_25_21, output_MAC_25_22, output_MAC_25_23, output_MAC_25_24, output_MAC_25_25, output_MAC_25_26, output_MAC_25_27, output_MAC_25_28, output_MAC_25_29, 
		output_MAC_25_30, output_MAC_25_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_26_0, output_MAC_26_1, output_MAC_26_2, output_MAC_26_3, output_MAC_26_4, output_MAC_26_5, output_MAC_26_6, output_MAC_26_7, output_MAC_26_8, output_MAC_26_9, 
		output_MAC_26_10, output_MAC_26_11, output_MAC_26_12, output_MAC_26_13, output_MAC_26_14, output_MAC_26_15, output_MAC_26_16, output_MAC_26_17, output_MAC_26_18, output_MAC_26_19, 
		output_MAC_26_20, output_MAC_26_21, output_MAC_26_22, output_MAC_26_23, output_MAC_26_24, output_MAC_26_25, output_MAC_26_26, output_MAC_26_27, output_MAC_26_28, output_MAC_26_29, 
		output_MAC_26_30, output_MAC_26_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_27_0, output_MAC_27_1, output_MAC_27_2, output_MAC_27_3, output_MAC_27_4, output_MAC_27_5, output_MAC_27_6, output_MAC_27_7, output_MAC_27_8, output_MAC_27_9, 
		output_MAC_27_10, output_MAC_27_11, output_MAC_27_12, output_MAC_27_13, output_MAC_27_14, output_MAC_27_15, output_MAC_27_16, output_MAC_27_17, output_MAC_27_18, output_MAC_27_19, 
		output_MAC_27_20, output_MAC_27_21, output_MAC_27_22, output_MAC_27_23, output_MAC_27_24, output_MAC_27_25, output_MAC_27_26, output_MAC_27_27, output_MAC_27_28, output_MAC_27_29, 
		output_MAC_27_30, output_MAC_27_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_28_0, output_MAC_28_1, output_MAC_28_2, output_MAC_28_3, output_MAC_28_4, output_MAC_28_5, output_MAC_28_6, output_MAC_28_7, output_MAC_28_8, output_MAC_28_9, 
		output_MAC_28_10, output_MAC_28_11, output_MAC_28_12, output_MAC_28_13, output_MAC_28_14, output_MAC_28_15, output_MAC_28_16, output_MAC_28_17, output_MAC_28_18, output_MAC_28_19, 
		output_MAC_28_20, output_MAC_28_21, output_MAC_28_22, output_MAC_28_23, output_MAC_28_24, output_MAC_28_25, output_MAC_28_26, output_MAC_28_27, output_MAC_28_28, output_MAC_28_29, 
		output_MAC_28_30, output_MAC_28_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_29_0, output_MAC_29_1, output_MAC_29_2, output_MAC_29_3, output_MAC_29_4, output_MAC_29_5, output_MAC_29_6, output_MAC_29_7, output_MAC_29_8, output_MAC_29_9, 
		output_MAC_29_10, output_MAC_29_11, output_MAC_29_12, output_MAC_29_13, output_MAC_29_14, output_MAC_29_15, output_MAC_29_16, output_MAC_29_17, output_MAC_29_18, output_MAC_29_19, 
		output_MAC_29_20, output_MAC_29_21, output_MAC_29_22, output_MAC_29_23, output_MAC_29_24, output_MAC_29_25, output_MAC_29_26, output_MAC_29_27, output_MAC_29_28, output_MAC_29_29, 
		output_MAC_29_30, output_MAC_29_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_30_0, output_MAC_30_1, output_MAC_30_2, output_MAC_30_3, output_MAC_30_4, output_MAC_30_5, output_MAC_30_6, output_MAC_30_7, output_MAC_30_8, output_MAC_30_9, 
		output_MAC_30_10, output_MAC_30_11, output_MAC_30_12, output_MAC_30_13, output_MAC_30_14, output_MAC_30_15, output_MAC_30_16, output_MAC_30_17, output_MAC_30_18, output_MAC_30_19, 
		output_MAC_30_20, output_MAC_30_21, output_MAC_30_22, output_MAC_30_23, output_MAC_30_24, output_MAC_30_25, output_MAC_30_26, output_MAC_30_27, output_MAC_30_28, output_MAC_30_29, 
		output_MAC_30_30, output_MAC_30_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_31_0, output_MAC_31_1, output_MAC_31_2, output_MAC_31_3, output_MAC_31_4, output_MAC_31_5, output_MAC_31_6, output_MAC_31_7, output_MAC_31_8, output_MAC_31_9, 
		output_MAC_31_10, output_MAC_31_11, output_MAC_31_12, output_MAC_31_13, output_MAC_31_14, output_MAC_31_15, output_MAC_31_16, output_MAC_31_17, output_MAC_31_18, output_MAC_31_19, 
		output_MAC_31_20, output_MAC_31_21, output_MAC_31_22, output_MAC_31_23, output_MAC_31_24, output_MAC_31_25, output_MAC_31_26, output_MAC_31_27, output_MAC_31_28, output_MAC_31_29, 
		output_MAC_31_30, output_MAC_31_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_32_0, output_MAC_32_1, output_MAC_32_2, output_MAC_32_3, output_MAC_32_4, output_MAC_32_5, output_MAC_32_6, output_MAC_32_7, output_MAC_32_8, output_MAC_32_9, 
		output_MAC_32_10, output_MAC_32_11, output_MAC_32_12, output_MAC_32_13, output_MAC_32_14, output_MAC_32_15, output_MAC_32_16, output_MAC_32_17, output_MAC_32_18, output_MAC_32_19, 
		output_MAC_32_20, output_MAC_32_21, output_MAC_32_22, output_MAC_32_23, output_MAC_32_24, output_MAC_32_25, output_MAC_32_26, output_MAC_32_27, output_MAC_32_28, output_MAC_32_29, 
		output_MAC_32_30, output_MAC_32_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_33_0, output_MAC_33_1, output_MAC_33_2, output_MAC_33_3, output_MAC_33_4, output_MAC_33_5, output_MAC_33_6, output_MAC_33_7, output_MAC_33_8, output_MAC_33_9, 
		output_MAC_33_10, output_MAC_33_11, output_MAC_33_12, output_MAC_33_13, output_MAC_33_14, output_MAC_33_15, output_MAC_33_16, output_MAC_33_17, output_MAC_33_18, output_MAC_33_19, 
		output_MAC_33_20, output_MAC_33_21, output_MAC_33_22, output_MAC_33_23, output_MAC_33_24, output_MAC_33_25, output_MAC_33_26, output_MAC_33_27, output_MAC_33_28, output_MAC_33_29, 
		output_MAC_33_30, output_MAC_33_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_34_0, output_MAC_34_1, output_MAC_34_2, output_MAC_34_3, output_MAC_34_4, output_MAC_34_5, output_MAC_34_6, output_MAC_34_7, output_MAC_34_8, output_MAC_34_9, 
		output_MAC_34_10, output_MAC_34_11, output_MAC_34_12, output_MAC_34_13, output_MAC_34_14, output_MAC_34_15, output_MAC_34_16, output_MAC_34_17, output_MAC_34_18, output_MAC_34_19, 
		output_MAC_34_20, output_MAC_34_21, output_MAC_34_22, output_MAC_34_23, output_MAC_34_24, output_MAC_34_25, output_MAC_34_26, output_MAC_34_27, output_MAC_34_28, output_MAC_34_29, 
		output_MAC_34_30, output_MAC_34_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_35_0, output_MAC_35_1, output_MAC_35_2, output_MAC_35_3, output_MAC_35_4, output_MAC_35_5, output_MAC_35_6, output_MAC_35_7, output_MAC_35_8, output_MAC_35_9, 
		output_MAC_35_10, output_MAC_35_11, output_MAC_35_12, output_MAC_35_13, output_MAC_35_14, output_MAC_35_15, output_MAC_35_16, output_MAC_35_17, output_MAC_35_18, output_MAC_35_19, 
		output_MAC_35_20, output_MAC_35_21, output_MAC_35_22, output_MAC_35_23, output_MAC_35_24, output_MAC_35_25, output_MAC_35_26, output_MAC_35_27, output_MAC_35_28, output_MAC_35_29, 
		output_MAC_35_30, output_MAC_35_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_36_0, output_MAC_36_1, output_MAC_36_2, output_MAC_36_3, output_MAC_36_4, output_MAC_36_5, output_MAC_36_6, output_MAC_36_7, output_MAC_36_8, output_MAC_36_9, 
		output_MAC_36_10, output_MAC_36_11, output_MAC_36_12, output_MAC_36_13, output_MAC_36_14, output_MAC_36_15, output_MAC_36_16, output_MAC_36_17, output_MAC_36_18, output_MAC_36_19, 
		output_MAC_36_20, output_MAC_36_21, output_MAC_36_22, output_MAC_36_23, output_MAC_36_24, output_MAC_36_25, output_MAC_36_26, output_MAC_36_27, output_MAC_36_28, output_MAC_36_29, 
		output_MAC_36_30, output_MAC_36_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_37_0, output_MAC_37_1, output_MAC_37_2, output_MAC_37_3, output_MAC_37_4, output_MAC_37_5, output_MAC_37_6, output_MAC_37_7, output_MAC_37_8, output_MAC_37_9, 
		output_MAC_37_10, output_MAC_37_11, output_MAC_37_12, output_MAC_37_13, output_MAC_37_14, output_MAC_37_15, output_MAC_37_16, output_MAC_37_17, output_MAC_37_18, output_MAC_37_19, 
		output_MAC_37_20, output_MAC_37_21, output_MAC_37_22, output_MAC_37_23, output_MAC_37_24, output_MAC_37_25, output_MAC_37_26, output_MAC_37_27, output_MAC_37_28, output_MAC_37_29, 
		output_MAC_37_30, output_MAC_37_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_38_0, output_MAC_38_1, output_MAC_38_2, output_MAC_38_3, output_MAC_38_4, output_MAC_38_5, output_MAC_38_6, output_MAC_38_7, output_MAC_38_8, output_MAC_38_9, 
		output_MAC_38_10, output_MAC_38_11, output_MAC_38_12, output_MAC_38_13, output_MAC_38_14, output_MAC_38_15, output_MAC_38_16, output_MAC_38_17, output_MAC_38_18, output_MAC_38_19, 
		output_MAC_38_20, output_MAC_38_21, output_MAC_38_22, output_MAC_38_23, output_MAC_38_24, output_MAC_38_25, output_MAC_38_26, output_MAC_38_27, output_MAC_38_28, output_MAC_38_29, 
		output_MAC_38_30, output_MAC_38_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_39_0, output_MAC_39_1, output_MAC_39_2, output_MAC_39_3, output_MAC_39_4, output_MAC_39_5, output_MAC_39_6, output_MAC_39_7, output_MAC_39_8, output_MAC_39_9, 
		output_MAC_39_10, output_MAC_39_11, output_MAC_39_12, output_MAC_39_13, output_MAC_39_14, output_MAC_39_15, output_MAC_39_16, output_MAC_39_17, output_MAC_39_18, output_MAC_39_19, 
		output_MAC_39_20, output_MAC_39_21, output_MAC_39_22, output_MAC_39_23, output_MAC_39_24, output_MAC_39_25, output_MAC_39_26, output_MAC_39_27, output_MAC_39_28, output_MAC_39_29, 
		output_MAC_39_30, output_MAC_39_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_40_0, output_MAC_40_1, output_MAC_40_2, output_MAC_40_3, output_MAC_40_4, output_MAC_40_5, output_MAC_40_6, output_MAC_40_7, output_MAC_40_8, output_MAC_40_9, 
		output_MAC_40_10, output_MAC_40_11, output_MAC_40_12, output_MAC_40_13, output_MAC_40_14, output_MAC_40_15, output_MAC_40_16, output_MAC_40_17, output_MAC_40_18, output_MAC_40_19, 
		output_MAC_40_20, output_MAC_40_21, output_MAC_40_22, output_MAC_40_23, output_MAC_40_24, output_MAC_40_25, output_MAC_40_26, output_MAC_40_27, output_MAC_40_28, output_MAC_40_29, 
		output_MAC_40_30, output_MAC_40_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_41_0, output_MAC_41_1, output_MAC_41_2, output_MAC_41_3, output_MAC_41_4, output_MAC_41_5, output_MAC_41_6, output_MAC_41_7, output_MAC_41_8, output_MAC_41_9, 
		output_MAC_41_10, output_MAC_41_11, output_MAC_41_12, output_MAC_41_13, output_MAC_41_14, output_MAC_41_15, output_MAC_41_16, output_MAC_41_17, output_MAC_41_18, output_MAC_41_19, 
		output_MAC_41_20, output_MAC_41_21, output_MAC_41_22, output_MAC_41_23, output_MAC_41_24, output_MAC_41_25, output_MAC_41_26, output_MAC_41_27, output_MAC_41_28, output_MAC_41_29, 
		output_MAC_41_30, output_MAC_41_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_42_0, output_MAC_42_1, output_MAC_42_2, output_MAC_42_3, output_MAC_42_4, output_MAC_42_5, output_MAC_42_6, output_MAC_42_7, output_MAC_42_8, output_MAC_42_9, 
		output_MAC_42_10, output_MAC_42_11, output_MAC_42_12, output_MAC_42_13, output_MAC_42_14, output_MAC_42_15, output_MAC_42_16, output_MAC_42_17, output_MAC_42_18, output_MAC_42_19, 
		output_MAC_42_20, output_MAC_42_21, output_MAC_42_22, output_MAC_42_23, output_MAC_42_24, output_MAC_42_25, output_MAC_42_26, output_MAC_42_27, output_MAC_42_28, output_MAC_42_29, 
		output_MAC_42_30, output_MAC_42_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_43_0, output_MAC_43_1, output_MAC_43_2, output_MAC_43_3, output_MAC_43_4, output_MAC_43_5, output_MAC_43_6, output_MAC_43_7, output_MAC_43_8, output_MAC_43_9, 
		output_MAC_43_10, output_MAC_43_11, output_MAC_43_12, output_MAC_43_13, output_MAC_43_14, output_MAC_43_15, output_MAC_43_16, output_MAC_43_17, output_MAC_43_18, output_MAC_43_19, 
		output_MAC_43_20, output_MAC_43_21, output_MAC_43_22, output_MAC_43_23, output_MAC_43_24, output_MAC_43_25, output_MAC_43_26, output_MAC_43_27, output_MAC_43_28, output_MAC_43_29, 
		output_MAC_43_30, output_MAC_43_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_44_0, output_MAC_44_1, output_MAC_44_2, output_MAC_44_3, output_MAC_44_4, output_MAC_44_5, output_MAC_44_6, output_MAC_44_7, output_MAC_44_8, output_MAC_44_9, 
		output_MAC_44_10, output_MAC_44_11, output_MAC_44_12, output_MAC_44_13, output_MAC_44_14, output_MAC_44_15, output_MAC_44_16, output_MAC_44_17, output_MAC_44_18, output_MAC_44_19, 
		output_MAC_44_20, output_MAC_44_21, output_MAC_44_22, output_MAC_44_23, output_MAC_44_24, output_MAC_44_25, output_MAC_44_26, output_MAC_44_27, output_MAC_44_28, output_MAC_44_29, 
		output_MAC_44_30, output_MAC_44_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_45_0, output_MAC_45_1, output_MAC_45_2, output_MAC_45_3, output_MAC_45_4, output_MAC_45_5, output_MAC_45_6, output_MAC_45_7, output_MAC_45_8, output_MAC_45_9, 
		output_MAC_45_10, output_MAC_45_11, output_MAC_45_12, output_MAC_45_13, output_MAC_45_14, output_MAC_45_15, output_MAC_45_16, output_MAC_45_17, output_MAC_45_18, output_MAC_45_19, 
		output_MAC_45_20, output_MAC_45_21, output_MAC_45_22, output_MAC_45_23, output_MAC_45_24, output_MAC_45_25, output_MAC_45_26, output_MAC_45_27, output_MAC_45_28, output_MAC_45_29, 
		output_MAC_45_30, output_MAC_45_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_46_0, output_MAC_46_1, output_MAC_46_2, output_MAC_46_3, output_MAC_46_4, output_MAC_46_5, output_MAC_46_6, output_MAC_46_7, output_MAC_46_8, output_MAC_46_9, 
		output_MAC_46_10, output_MAC_46_11, output_MAC_46_12, output_MAC_46_13, output_MAC_46_14, output_MAC_46_15, output_MAC_46_16, output_MAC_46_17, output_MAC_46_18, output_MAC_46_19, 
		output_MAC_46_20, output_MAC_46_21, output_MAC_46_22, output_MAC_46_23, output_MAC_46_24, output_MAC_46_25, output_MAC_46_26, output_MAC_46_27, output_MAC_46_28, output_MAC_46_29, 
		output_MAC_46_30, output_MAC_46_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_47_0, output_MAC_47_1, output_MAC_47_2, output_MAC_47_3, output_MAC_47_4, output_MAC_47_5, output_MAC_47_6, output_MAC_47_7, output_MAC_47_8, output_MAC_47_9, 
		output_MAC_47_10, output_MAC_47_11, output_MAC_47_12, output_MAC_47_13, output_MAC_47_14, output_MAC_47_15, output_MAC_47_16, output_MAC_47_17, output_MAC_47_18, output_MAC_47_19, 
		output_MAC_47_20, output_MAC_47_21, output_MAC_47_22, output_MAC_47_23, output_MAC_47_24, output_MAC_47_25, output_MAC_47_26, output_MAC_47_27, output_MAC_47_28, output_MAC_47_29, 
		output_MAC_47_30, output_MAC_47_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_48_0, output_MAC_48_1, output_MAC_48_2, output_MAC_48_3, output_MAC_48_4, output_MAC_48_5, output_MAC_48_6, output_MAC_48_7, output_MAC_48_8, output_MAC_48_9, 
		output_MAC_48_10, output_MAC_48_11, output_MAC_48_12, output_MAC_48_13, output_MAC_48_14, output_MAC_48_15, output_MAC_48_16, output_MAC_48_17, output_MAC_48_18, output_MAC_48_19, 
		output_MAC_48_20, output_MAC_48_21, output_MAC_48_22, output_MAC_48_23, output_MAC_48_24, output_MAC_48_25, output_MAC_48_26, output_MAC_48_27, output_MAC_48_28, output_MAC_48_29, 
		output_MAC_48_30, output_MAC_48_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_49_0, output_MAC_49_1, output_MAC_49_2, output_MAC_49_3, output_MAC_49_4, output_MAC_49_5, output_MAC_49_6, output_MAC_49_7, output_MAC_49_8, output_MAC_49_9, 
		output_MAC_49_10, output_MAC_49_11, output_MAC_49_12, output_MAC_49_13, output_MAC_49_14, output_MAC_49_15, output_MAC_49_16, output_MAC_49_17, output_MAC_49_18, output_MAC_49_19, 
		output_MAC_49_20, output_MAC_49_21, output_MAC_49_22, output_MAC_49_23, output_MAC_49_24, output_MAC_49_25, output_MAC_49_26, output_MAC_49_27, output_MAC_49_28, output_MAC_49_29, 
		output_MAC_49_30, output_MAC_49_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_50_0, output_MAC_50_1, output_MAC_50_2, output_MAC_50_3, output_MAC_50_4, output_MAC_50_5, output_MAC_50_6, output_MAC_50_7, output_MAC_50_8, output_MAC_50_9, 
		output_MAC_50_10, output_MAC_50_11, output_MAC_50_12, output_MAC_50_13, output_MAC_50_14, output_MAC_50_15, output_MAC_50_16, output_MAC_50_17, output_MAC_50_18, output_MAC_50_19, 
		output_MAC_50_20, output_MAC_50_21, output_MAC_50_22, output_MAC_50_23, output_MAC_50_24, output_MAC_50_25, output_MAC_50_26, output_MAC_50_27, output_MAC_50_28, output_MAC_50_29, 
		output_MAC_50_30, output_MAC_50_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_51_0, output_MAC_51_1, output_MAC_51_2, output_MAC_51_3, output_MAC_51_4, output_MAC_51_5, output_MAC_51_6, output_MAC_51_7, output_MAC_51_8, output_MAC_51_9, 
		output_MAC_51_10, output_MAC_51_11, output_MAC_51_12, output_MAC_51_13, output_MAC_51_14, output_MAC_51_15, output_MAC_51_16, output_MAC_51_17, output_MAC_51_18, output_MAC_51_19, 
		output_MAC_51_20, output_MAC_51_21, output_MAC_51_22, output_MAC_51_23, output_MAC_51_24, output_MAC_51_25, output_MAC_51_26, output_MAC_51_27, output_MAC_51_28, output_MAC_51_29, 
		output_MAC_51_30, output_MAC_51_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_52_0, output_MAC_52_1, output_MAC_52_2, output_MAC_52_3, output_MAC_52_4, output_MAC_52_5, output_MAC_52_6, output_MAC_52_7, output_MAC_52_8, output_MAC_52_9, 
		output_MAC_52_10, output_MAC_52_11, output_MAC_52_12, output_MAC_52_13, output_MAC_52_14, output_MAC_52_15, output_MAC_52_16, output_MAC_52_17, output_MAC_52_18, output_MAC_52_19, 
		output_MAC_52_20, output_MAC_52_21, output_MAC_52_22, output_MAC_52_23, output_MAC_52_24, output_MAC_52_25, output_MAC_52_26, output_MAC_52_27, output_MAC_52_28, output_MAC_52_29, 
		output_MAC_52_30, output_MAC_52_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_53_0, output_MAC_53_1, output_MAC_53_2, output_MAC_53_3, output_MAC_53_4, output_MAC_53_5, output_MAC_53_6, output_MAC_53_7, output_MAC_53_8, output_MAC_53_9, 
		output_MAC_53_10, output_MAC_53_11, output_MAC_53_12, output_MAC_53_13, output_MAC_53_14, output_MAC_53_15, output_MAC_53_16, output_MAC_53_17, output_MAC_53_18, output_MAC_53_19, 
		output_MAC_53_20, output_MAC_53_21, output_MAC_53_22, output_MAC_53_23, output_MAC_53_24, output_MAC_53_25, output_MAC_53_26, output_MAC_53_27, output_MAC_53_28, output_MAC_53_29, 
		output_MAC_53_30, output_MAC_53_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_54_0, output_MAC_54_1, output_MAC_54_2, output_MAC_54_3, output_MAC_54_4, output_MAC_54_5, output_MAC_54_6, output_MAC_54_7, output_MAC_54_8, output_MAC_54_9, 
		output_MAC_54_10, output_MAC_54_11, output_MAC_54_12, output_MAC_54_13, output_MAC_54_14, output_MAC_54_15, output_MAC_54_16, output_MAC_54_17, output_MAC_54_18, output_MAC_54_19, 
		output_MAC_54_20, output_MAC_54_21, output_MAC_54_22, output_MAC_54_23, output_MAC_54_24, output_MAC_54_25, output_MAC_54_26, output_MAC_54_27, output_MAC_54_28, output_MAC_54_29, 
		output_MAC_54_30, output_MAC_54_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_55_0, output_MAC_55_1, output_MAC_55_2, output_MAC_55_3, output_MAC_55_4, output_MAC_55_5, output_MAC_55_6, output_MAC_55_7, output_MAC_55_8, output_MAC_55_9, 
		output_MAC_55_10, output_MAC_55_11, output_MAC_55_12, output_MAC_55_13, output_MAC_55_14, output_MAC_55_15, output_MAC_55_16, output_MAC_55_17, output_MAC_55_18, output_MAC_55_19, 
		output_MAC_55_20, output_MAC_55_21, output_MAC_55_22, output_MAC_55_23, output_MAC_55_24, output_MAC_55_25, output_MAC_55_26, output_MAC_55_27, output_MAC_55_28, output_MAC_55_29, 
		output_MAC_55_30, output_MAC_55_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_56_0, output_MAC_56_1, output_MAC_56_2, output_MAC_56_3, output_MAC_56_4, output_MAC_56_5, output_MAC_56_6, output_MAC_56_7, output_MAC_56_8, output_MAC_56_9, 
		output_MAC_56_10, output_MAC_56_11, output_MAC_56_12, output_MAC_56_13, output_MAC_56_14, output_MAC_56_15, output_MAC_56_16, output_MAC_56_17, output_MAC_56_18, output_MAC_56_19, 
		output_MAC_56_20, output_MAC_56_21, output_MAC_56_22, output_MAC_56_23, output_MAC_56_24, output_MAC_56_25, output_MAC_56_26, output_MAC_56_27, output_MAC_56_28, output_MAC_56_29, 
		output_MAC_56_30, output_MAC_56_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_57_0, output_MAC_57_1, output_MAC_57_2, output_MAC_57_3, output_MAC_57_4, output_MAC_57_5, output_MAC_57_6, output_MAC_57_7, output_MAC_57_8, output_MAC_57_9, 
		output_MAC_57_10, output_MAC_57_11, output_MAC_57_12, output_MAC_57_13, output_MAC_57_14, output_MAC_57_15, output_MAC_57_16, output_MAC_57_17, output_MAC_57_18, output_MAC_57_19, 
		output_MAC_57_20, output_MAC_57_21, output_MAC_57_22, output_MAC_57_23, output_MAC_57_24, output_MAC_57_25, output_MAC_57_26, output_MAC_57_27, output_MAC_57_28, output_MAC_57_29, 
		output_MAC_57_30, output_MAC_57_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_58_0, output_MAC_58_1, output_MAC_58_2, output_MAC_58_3, output_MAC_58_4, output_MAC_58_5, output_MAC_58_6, output_MAC_58_7, output_MAC_58_8, output_MAC_58_9, 
		output_MAC_58_10, output_MAC_58_11, output_MAC_58_12, output_MAC_58_13, output_MAC_58_14, output_MAC_58_15, output_MAC_58_16, output_MAC_58_17, output_MAC_58_18, output_MAC_58_19, 
		output_MAC_58_20, output_MAC_58_21, output_MAC_58_22, output_MAC_58_23, output_MAC_58_24, output_MAC_58_25, output_MAC_58_26, output_MAC_58_27, output_MAC_58_28, output_MAC_58_29, 
		output_MAC_58_30, output_MAC_58_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_59_0, output_MAC_59_1, output_MAC_59_2, output_MAC_59_3, output_MAC_59_4, output_MAC_59_5, output_MAC_59_6, output_MAC_59_7, output_MAC_59_8, output_MAC_59_9, 
		output_MAC_59_10, output_MAC_59_11, output_MAC_59_12, output_MAC_59_13, output_MAC_59_14, output_MAC_59_15, output_MAC_59_16, output_MAC_59_17, output_MAC_59_18, output_MAC_59_19, 
		output_MAC_59_20, output_MAC_59_21, output_MAC_59_22, output_MAC_59_23, output_MAC_59_24, output_MAC_59_25, output_MAC_59_26, output_MAC_59_27, output_MAC_59_28, output_MAC_59_29, 
		output_MAC_59_30, output_MAC_59_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_60_0, output_MAC_60_1, output_MAC_60_2, output_MAC_60_3, output_MAC_60_4, output_MAC_60_5, output_MAC_60_6, output_MAC_60_7, output_MAC_60_8, output_MAC_60_9, 
		output_MAC_60_10, output_MAC_60_11, output_MAC_60_12, output_MAC_60_13, output_MAC_60_14, output_MAC_60_15, output_MAC_60_16, output_MAC_60_17, output_MAC_60_18, output_MAC_60_19, 
		output_MAC_60_20, output_MAC_60_21, output_MAC_60_22, output_MAC_60_23, output_MAC_60_24, output_MAC_60_25, output_MAC_60_26, output_MAC_60_27, output_MAC_60_28, output_MAC_60_29, 
		output_MAC_60_30, output_MAC_60_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_61_0, output_MAC_61_1, output_MAC_61_2, output_MAC_61_3, output_MAC_61_4, output_MAC_61_5, output_MAC_61_6, output_MAC_61_7, output_MAC_61_8, output_MAC_61_9, 
		output_MAC_61_10, output_MAC_61_11, output_MAC_61_12, output_MAC_61_13, output_MAC_61_14, output_MAC_61_15, output_MAC_61_16, output_MAC_61_17, output_MAC_61_18, output_MAC_61_19, 
		output_MAC_61_20, output_MAC_61_21, output_MAC_61_22, output_MAC_61_23, output_MAC_61_24, output_MAC_61_25, output_MAC_61_26, output_MAC_61_27, output_MAC_61_28, output_MAC_61_29, 
		output_MAC_61_30, output_MAC_61_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_62_0, output_MAC_62_1, output_MAC_62_2, output_MAC_62_3, output_MAC_62_4, output_MAC_62_5, output_MAC_62_6, output_MAC_62_7, output_MAC_62_8, output_MAC_62_9, 
		output_MAC_62_10, output_MAC_62_11, output_MAC_62_12, output_MAC_62_13, output_MAC_62_14, output_MAC_62_15, output_MAC_62_16, output_MAC_62_17, output_MAC_62_18, output_MAC_62_19, 
		output_MAC_62_20, output_MAC_62_21, output_MAC_62_22, output_MAC_62_23, output_MAC_62_24, output_MAC_62_25, output_MAC_62_26, output_MAC_62_27, output_MAC_62_28, output_MAC_62_29, 
		output_MAC_62_30, output_MAC_62_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_63_0, output_MAC_63_1, output_MAC_63_2, output_MAC_63_3, output_MAC_63_4, output_MAC_63_5, output_MAC_63_6, output_MAC_63_7, output_MAC_63_8, output_MAC_63_9, 
		output_MAC_63_10, output_MAC_63_11, output_MAC_63_12, output_MAC_63_13, output_MAC_63_14, output_MAC_63_15, output_MAC_63_16, output_MAC_63_17, output_MAC_63_18, output_MAC_63_19, 
		output_MAC_63_20, output_MAC_63_21, output_MAC_63_22, output_MAC_63_23, output_MAC_63_24, output_MAC_63_25, output_MAC_63_26, output_MAC_63_27, output_MAC_63_28, output_MAC_63_29, 
		output_MAC_63_30, output_MAC_63_31: STD_LOGIC_VECTOR(31 downto 0);

BEGIN

	MAC_0_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_0, data_out=>output_MAC_0_0);
	MAC_0_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_1, data_out=>output_MAC_0_1);
	MAC_0_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_2, data_out=>output_MAC_0_2);
	MAC_0_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_3, data_out=>output_MAC_0_3);
	MAC_0_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_4, data_out=>output_MAC_0_4);
	MAC_0_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_5, data_out=>output_MAC_0_5);
	MAC_0_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_6, data_out=>output_MAC_0_6);
	MAC_0_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_7, data_out=>output_MAC_0_7);
	MAC_0_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_8, data_out=>output_MAC_0_8);
	MAC_0_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_9, data_out=>output_MAC_0_9);
	MAC_0_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_10, data_out=>output_MAC_0_10);
	MAC_0_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_11, data_out=>output_MAC_0_11);
	MAC_0_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_12, data_out=>output_MAC_0_12);
	MAC_0_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_13, data_out=>output_MAC_0_13);
	MAC_0_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_14, data_out=>output_MAC_0_14);
	MAC_0_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_15, data_out=>output_MAC_0_15);
	MAC_0_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_16, data_out=>output_MAC_0_16);
	MAC_0_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_17, data_out=>output_MAC_0_17);
	MAC_0_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_18, data_out=>output_MAC_0_18);
	MAC_0_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_19, data_out=>output_MAC_0_19);
	MAC_0_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_20, data_out=>output_MAC_0_20);
	MAC_0_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_21, data_out=>output_MAC_0_21);
	MAC_0_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_22, data_out=>output_MAC_0_22);
	MAC_0_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_23, data_out=>output_MAC_0_23);
	MAC_0_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_24, data_out=>output_MAC_0_24);
	MAC_0_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_25, data_out=>output_MAC_0_25);
	MAC_0_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_26, data_out=>output_MAC_0_26);
	MAC_0_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_27, data_out=>output_MAC_0_27);
	MAC_0_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_28, data_out=>output_MAC_0_28);
	MAC_0_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_29, data_out=>output_MAC_0_29);
	MAC_0_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_30, data_out=>output_MAC_0_30);
	MAC_0_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_31, data_out=>output_MAC_0_31);
	MAC_1_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_0, data_out=>output_MAC_1_0);
	MAC_1_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_1, data_out=>output_MAC_1_1);
	MAC_1_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_2, data_out=>output_MAC_1_2);
	MAC_1_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_3, data_out=>output_MAC_1_3);
	MAC_1_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_4, data_out=>output_MAC_1_4);
	MAC_1_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_5, data_out=>output_MAC_1_5);
	MAC_1_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_6, data_out=>output_MAC_1_6);
	MAC_1_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_7, data_out=>output_MAC_1_7);
	MAC_1_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_8, data_out=>output_MAC_1_8);
	MAC_1_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_9, data_out=>output_MAC_1_9);
	MAC_1_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_10, data_out=>output_MAC_1_10);
	MAC_1_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_11, data_out=>output_MAC_1_11);
	MAC_1_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_12, data_out=>output_MAC_1_12);
	MAC_1_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_13, data_out=>output_MAC_1_13);
	MAC_1_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_14, data_out=>output_MAC_1_14);
	MAC_1_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_15, data_out=>output_MAC_1_15);
	MAC_1_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_16, data_out=>output_MAC_1_16);
	MAC_1_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_17, data_out=>output_MAC_1_17);
	MAC_1_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_18, data_out=>output_MAC_1_18);
	MAC_1_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_19, data_out=>output_MAC_1_19);
	MAC_1_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_20, data_out=>output_MAC_1_20);
	MAC_1_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_21, data_out=>output_MAC_1_21);
	MAC_1_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_22, data_out=>output_MAC_1_22);
	MAC_1_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_23, data_out=>output_MAC_1_23);
	MAC_1_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_24, data_out=>output_MAC_1_24);
	MAC_1_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_25, data_out=>output_MAC_1_25);
	MAC_1_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_26, data_out=>output_MAC_1_26);
	MAC_1_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_27, data_out=>output_MAC_1_27);
	MAC_1_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_28, data_out=>output_MAC_1_28);
	MAC_1_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_29, data_out=>output_MAC_1_29);
	MAC_1_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_30, data_out=>output_MAC_1_30);
	MAC_1_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_31, data_out=>output_MAC_1_31);
	MAC_2_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_0, data_out=>output_MAC_2_0);
	MAC_2_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_1, data_out=>output_MAC_2_1);
	MAC_2_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_2, data_out=>output_MAC_2_2);
	MAC_2_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_3, data_out=>output_MAC_2_3);
	MAC_2_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_4, data_out=>output_MAC_2_4);
	MAC_2_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_5, data_out=>output_MAC_2_5);
	MAC_2_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_6, data_out=>output_MAC_2_6);
	MAC_2_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_7, data_out=>output_MAC_2_7);
	MAC_2_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_8, data_out=>output_MAC_2_8);
	MAC_2_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_9, data_out=>output_MAC_2_9);
	MAC_2_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_10, data_out=>output_MAC_2_10);
	MAC_2_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_11, data_out=>output_MAC_2_11);
	MAC_2_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_12, data_out=>output_MAC_2_12);
	MAC_2_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_13, data_out=>output_MAC_2_13);
	MAC_2_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_14, data_out=>output_MAC_2_14);
	MAC_2_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_15, data_out=>output_MAC_2_15);
	MAC_2_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_16, data_out=>output_MAC_2_16);
	MAC_2_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_17, data_out=>output_MAC_2_17);
	MAC_2_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_18, data_out=>output_MAC_2_18);
	MAC_2_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_19, data_out=>output_MAC_2_19);
	MAC_2_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_20, data_out=>output_MAC_2_20);
	MAC_2_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_21, data_out=>output_MAC_2_21);
	MAC_2_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_22, data_out=>output_MAC_2_22);
	MAC_2_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_23, data_out=>output_MAC_2_23);
	MAC_2_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_24, data_out=>output_MAC_2_24);
	MAC_2_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_25, data_out=>output_MAC_2_25);
	MAC_2_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_26, data_out=>output_MAC_2_26);
	MAC_2_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_27, data_out=>output_MAC_2_27);
	MAC_2_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_28, data_out=>output_MAC_2_28);
	MAC_2_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_29, data_out=>output_MAC_2_29);
	MAC_2_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_30, data_out=>output_MAC_2_30);
	MAC_2_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_31, data_out=>output_MAC_2_31);
	MAC_3_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_0, data_out=>output_MAC_3_0);
	MAC_3_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_1, data_out=>output_MAC_3_1);
	MAC_3_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_2, data_out=>output_MAC_3_2);
	MAC_3_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_3, data_out=>output_MAC_3_3);
	MAC_3_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_4, data_out=>output_MAC_3_4);
	MAC_3_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_5, data_out=>output_MAC_3_5);
	MAC_3_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_6, data_out=>output_MAC_3_6);
	MAC_3_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_7, data_out=>output_MAC_3_7);
	MAC_3_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_8, data_out=>output_MAC_3_8);
	MAC_3_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_9, data_out=>output_MAC_3_9);
	MAC_3_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_10, data_out=>output_MAC_3_10);
	MAC_3_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_11, data_out=>output_MAC_3_11);
	MAC_3_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_12, data_out=>output_MAC_3_12);
	MAC_3_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_13, data_out=>output_MAC_3_13);
	MAC_3_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_14, data_out=>output_MAC_3_14);
	MAC_3_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_15, data_out=>output_MAC_3_15);
	MAC_3_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_16, data_out=>output_MAC_3_16);
	MAC_3_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_17, data_out=>output_MAC_3_17);
	MAC_3_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_18, data_out=>output_MAC_3_18);
	MAC_3_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_19, data_out=>output_MAC_3_19);
	MAC_3_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_20, data_out=>output_MAC_3_20);
	MAC_3_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_21, data_out=>output_MAC_3_21);
	MAC_3_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_22, data_out=>output_MAC_3_22);
	MAC_3_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_23, data_out=>output_MAC_3_23);
	MAC_3_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_24, data_out=>output_MAC_3_24);
	MAC_3_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_25, data_out=>output_MAC_3_25);
	MAC_3_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_26, data_out=>output_MAC_3_26);
	MAC_3_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_27, data_out=>output_MAC_3_27);
	MAC_3_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_28, data_out=>output_MAC_3_28);
	MAC_3_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_29, data_out=>output_MAC_3_29);
	MAC_3_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_30, data_out=>output_MAC_3_30);
	MAC_3_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_31, data_out=>output_MAC_3_31);
	MAC_4_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_0, data_out=>output_MAC_4_0);
	MAC_4_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_1, data_out=>output_MAC_4_1);
	MAC_4_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_2, data_out=>output_MAC_4_2);
	MAC_4_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_3, data_out=>output_MAC_4_3);
	MAC_4_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_4, data_out=>output_MAC_4_4);
	MAC_4_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_5, data_out=>output_MAC_4_5);
	MAC_4_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_6, data_out=>output_MAC_4_6);
	MAC_4_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_7, data_out=>output_MAC_4_7);
	MAC_4_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_8, data_out=>output_MAC_4_8);
	MAC_4_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_9, data_out=>output_MAC_4_9);
	MAC_4_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_10, data_out=>output_MAC_4_10);
	MAC_4_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_11, data_out=>output_MAC_4_11);
	MAC_4_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_12, data_out=>output_MAC_4_12);
	MAC_4_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_13, data_out=>output_MAC_4_13);
	MAC_4_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_14, data_out=>output_MAC_4_14);
	MAC_4_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_15, data_out=>output_MAC_4_15);
	MAC_4_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_16, data_out=>output_MAC_4_16);
	MAC_4_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_17, data_out=>output_MAC_4_17);
	MAC_4_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_18, data_out=>output_MAC_4_18);
	MAC_4_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_19, data_out=>output_MAC_4_19);
	MAC_4_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_20, data_out=>output_MAC_4_20);
	MAC_4_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_21, data_out=>output_MAC_4_21);
	MAC_4_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_22, data_out=>output_MAC_4_22);
	MAC_4_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_23, data_out=>output_MAC_4_23);
	MAC_4_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_24, data_out=>output_MAC_4_24);
	MAC_4_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_25, data_out=>output_MAC_4_25);
	MAC_4_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_26, data_out=>output_MAC_4_26);
	MAC_4_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_27, data_out=>output_MAC_4_27);
	MAC_4_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_28, data_out=>output_MAC_4_28);
	MAC_4_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_29, data_out=>output_MAC_4_29);
	MAC_4_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_30, data_out=>output_MAC_4_30);
	MAC_4_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_31, data_out=>output_MAC_4_31);
	MAC_5_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_0, data_out=>output_MAC_5_0);
	MAC_5_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_1, data_out=>output_MAC_5_1);
	MAC_5_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_2, data_out=>output_MAC_5_2);
	MAC_5_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_3, data_out=>output_MAC_5_3);
	MAC_5_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_4, data_out=>output_MAC_5_4);
	MAC_5_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_5, data_out=>output_MAC_5_5);
	MAC_5_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_6, data_out=>output_MAC_5_6);
	MAC_5_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_7, data_out=>output_MAC_5_7);
	MAC_5_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_8, data_out=>output_MAC_5_8);
	MAC_5_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_9, data_out=>output_MAC_5_9);
	MAC_5_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_10, data_out=>output_MAC_5_10);
	MAC_5_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_11, data_out=>output_MAC_5_11);
	MAC_5_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_12, data_out=>output_MAC_5_12);
	MAC_5_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_13, data_out=>output_MAC_5_13);
	MAC_5_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_14, data_out=>output_MAC_5_14);
	MAC_5_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_15, data_out=>output_MAC_5_15);
	MAC_5_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_16, data_out=>output_MAC_5_16);
	MAC_5_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_17, data_out=>output_MAC_5_17);
	MAC_5_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_18, data_out=>output_MAC_5_18);
	MAC_5_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_19, data_out=>output_MAC_5_19);
	MAC_5_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_20, data_out=>output_MAC_5_20);
	MAC_5_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_21, data_out=>output_MAC_5_21);
	MAC_5_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_22, data_out=>output_MAC_5_22);
	MAC_5_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_23, data_out=>output_MAC_5_23);
	MAC_5_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_24, data_out=>output_MAC_5_24);
	MAC_5_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_25, data_out=>output_MAC_5_25);
	MAC_5_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_26, data_out=>output_MAC_5_26);
	MAC_5_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_27, data_out=>output_MAC_5_27);
	MAC_5_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_28, data_out=>output_MAC_5_28);
	MAC_5_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_29, data_out=>output_MAC_5_29);
	MAC_5_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_30, data_out=>output_MAC_5_30);
	MAC_5_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_31, data_out=>output_MAC_5_31);
	MAC_6_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_0, data_out=>output_MAC_6_0);
	MAC_6_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_1, data_out=>output_MAC_6_1);
	MAC_6_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_2, data_out=>output_MAC_6_2);
	MAC_6_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_3, data_out=>output_MAC_6_3);
	MAC_6_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_4, data_out=>output_MAC_6_4);
	MAC_6_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_5, data_out=>output_MAC_6_5);
	MAC_6_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_6, data_out=>output_MAC_6_6);
	MAC_6_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_7, data_out=>output_MAC_6_7);
	MAC_6_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_8, data_out=>output_MAC_6_8);
	MAC_6_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_9, data_out=>output_MAC_6_9);
	MAC_6_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_10, data_out=>output_MAC_6_10);
	MAC_6_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_11, data_out=>output_MAC_6_11);
	MAC_6_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_12, data_out=>output_MAC_6_12);
	MAC_6_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_13, data_out=>output_MAC_6_13);
	MAC_6_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_14, data_out=>output_MAC_6_14);
	MAC_6_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_15, data_out=>output_MAC_6_15);
	MAC_6_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_16, data_out=>output_MAC_6_16);
	MAC_6_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_17, data_out=>output_MAC_6_17);
	MAC_6_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_18, data_out=>output_MAC_6_18);
	MAC_6_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_19, data_out=>output_MAC_6_19);
	MAC_6_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_20, data_out=>output_MAC_6_20);
	MAC_6_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_21, data_out=>output_MAC_6_21);
	MAC_6_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_22, data_out=>output_MAC_6_22);
	MAC_6_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_23, data_out=>output_MAC_6_23);
	MAC_6_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_24, data_out=>output_MAC_6_24);
	MAC_6_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_25, data_out=>output_MAC_6_25);
	MAC_6_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_26, data_out=>output_MAC_6_26);
	MAC_6_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_27, data_out=>output_MAC_6_27);
	MAC_6_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_28, data_out=>output_MAC_6_28);
	MAC_6_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_29, data_out=>output_MAC_6_29);
	MAC_6_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_30, data_out=>output_MAC_6_30);
	MAC_6_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_31, data_out=>output_MAC_6_31);
	MAC_7_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_0, data_out=>output_MAC_7_0);
	MAC_7_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_1, data_out=>output_MAC_7_1);
	MAC_7_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_2, data_out=>output_MAC_7_2);
	MAC_7_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_3, data_out=>output_MAC_7_3);
	MAC_7_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_4, data_out=>output_MAC_7_4);
	MAC_7_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_5, data_out=>output_MAC_7_5);
	MAC_7_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_6, data_out=>output_MAC_7_6);
	MAC_7_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_7, data_out=>output_MAC_7_7);
	MAC_7_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_8, data_out=>output_MAC_7_8);
	MAC_7_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_9, data_out=>output_MAC_7_9);
	MAC_7_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_10, data_out=>output_MAC_7_10);
	MAC_7_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_11, data_out=>output_MAC_7_11);
	MAC_7_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_12, data_out=>output_MAC_7_12);
	MAC_7_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_13, data_out=>output_MAC_7_13);
	MAC_7_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_14, data_out=>output_MAC_7_14);
	MAC_7_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_15, data_out=>output_MAC_7_15);
	MAC_7_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_16, data_out=>output_MAC_7_16);
	MAC_7_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_17, data_out=>output_MAC_7_17);
	MAC_7_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_18, data_out=>output_MAC_7_18);
	MAC_7_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_19, data_out=>output_MAC_7_19);
	MAC_7_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_20, data_out=>output_MAC_7_20);
	MAC_7_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_21, data_out=>output_MAC_7_21);
	MAC_7_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_22, data_out=>output_MAC_7_22);
	MAC_7_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_23, data_out=>output_MAC_7_23);
	MAC_7_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_24, data_out=>output_MAC_7_24);
	MAC_7_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_25, data_out=>output_MAC_7_25);
	MAC_7_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_26, data_out=>output_MAC_7_26);
	MAC_7_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_27, data_out=>output_MAC_7_27);
	MAC_7_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_28, data_out=>output_MAC_7_28);
	MAC_7_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_29, data_out=>output_MAC_7_29);
	MAC_7_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_30, data_out=>output_MAC_7_30);
	MAC_7_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_31, data_out=>output_MAC_7_31);
	MAC_8_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_0, data_out=>output_MAC_8_0);
	MAC_8_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_1, data_out=>output_MAC_8_1);
	MAC_8_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_2, data_out=>output_MAC_8_2);
	MAC_8_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_3, data_out=>output_MAC_8_3);
	MAC_8_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_4, data_out=>output_MAC_8_4);
	MAC_8_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_5, data_out=>output_MAC_8_5);
	MAC_8_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_6, data_out=>output_MAC_8_6);
	MAC_8_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_7, data_out=>output_MAC_8_7);
	MAC_8_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_8, data_out=>output_MAC_8_8);
	MAC_8_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_9, data_out=>output_MAC_8_9);
	MAC_8_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_10, data_out=>output_MAC_8_10);
	MAC_8_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_11, data_out=>output_MAC_8_11);
	MAC_8_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_12, data_out=>output_MAC_8_12);
	MAC_8_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_13, data_out=>output_MAC_8_13);
	MAC_8_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_14, data_out=>output_MAC_8_14);
	MAC_8_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_15, data_out=>output_MAC_8_15);
	MAC_8_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_16, data_out=>output_MAC_8_16);
	MAC_8_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_17, data_out=>output_MAC_8_17);
	MAC_8_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_18, data_out=>output_MAC_8_18);
	MAC_8_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_19, data_out=>output_MAC_8_19);
	MAC_8_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_20, data_out=>output_MAC_8_20);
	MAC_8_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_21, data_out=>output_MAC_8_21);
	MAC_8_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_22, data_out=>output_MAC_8_22);
	MAC_8_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_23, data_out=>output_MAC_8_23);
	MAC_8_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_24, data_out=>output_MAC_8_24);
	MAC_8_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_25, data_out=>output_MAC_8_25);
	MAC_8_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_26, data_out=>output_MAC_8_26);
	MAC_8_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_27, data_out=>output_MAC_8_27);
	MAC_8_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_28, data_out=>output_MAC_8_28);
	MAC_8_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_29, data_out=>output_MAC_8_29);
	MAC_8_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_30, data_out=>output_MAC_8_30);
	MAC_8_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_31, data_out=>output_MAC_8_31);
	MAC_9_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_0, data_out=>output_MAC_9_0);
	MAC_9_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_1, data_out=>output_MAC_9_1);
	MAC_9_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_2, data_out=>output_MAC_9_2);
	MAC_9_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_3, data_out=>output_MAC_9_3);
	MAC_9_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_4, data_out=>output_MAC_9_4);
	MAC_9_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_5, data_out=>output_MAC_9_5);
	MAC_9_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_6, data_out=>output_MAC_9_6);
	MAC_9_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_7, data_out=>output_MAC_9_7);
	MAC_9_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_8, data_out=>output_MAC_9_8);
	MAC_9_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_9, data_out=>output_MAC_9_9);
	MAC_9_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_10, data_out=>output_MAC_9_10);
	MAC_9_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_11, data_out=>output_MAC_9_11);
	MAC_9_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_12, data_out=>output_MAC_9_12);
	MAC_9_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_13, data_out=>output_MAC_9_13);
	MAC_9_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_14, data_out=>output_MAC_9_14);
	MAC_9_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_15, data_out=>output_MAC_9_15);
	MAC_9_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_16, data_out=>output_MAC_9_16);
	MAC_9_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_17, data_out=>output_MAC_9_17);
	MAC_9_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_18, data_out=>output_MAC_9_18);
	MAC_9_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_19, data_out=>output_MAC_9_19);
	MAC_9_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_20, data_out=>output_MAC_9_20);
	MAC_9_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_21, data_out=>output_MAC_9_21);
	MAC_9_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_22, data_out=>output_MAC_9_22);
	MAC_9_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_23, data_out=>output_MAC_9_23);
	MAC_9_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_24, data_out=>output_MAC_9_24);
	MAC_9_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_25, data_out=>output_MAC_9_25);
	MAC_9_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_26, data_out=>output_MAC_9_26);
	MAC_9_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_27, data_out=>output_MAC_9_27);
	MAC_9_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_28, data_out=>output_MAC_9_28);
	MAC_9_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_29, data_out=>output_MAC_9_29);
	MAC_9_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_30, data_out=>output_MAC_9_30);
	MAC_9_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_31, data_out=>output_MAC_9_31);
	MAC_10_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_0, data_out=>output_MAC_10_0);
	MAC_10_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_1, data_out=>output_MAC_10_1);
	MAC_10_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_2, data_out=>output_MAC_10_2);
	MAC_10_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_3, data_out=>output_MAC_10_3);
	MAC_10_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_4, data_out=>output_MAC_10_4);
	MAC_10_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_5, data_out=>output_MAC_10_5);
	MAC_10_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_6, data_out=>output_MAC_10_6);
	MAC_10_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_7, data_out=>output_MAC_10_7);
	MAC_10_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_8, data_out=>output_MAC_10_8);
	MAC_10_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_9, data_out=>output_MAC_10_9);
	MAC_10_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_10, data_out=>output_MAC_10_10);
	MAC_10_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_11, data_out=>output_MAC_10_11);
	MAC_10_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_12, data_out=>output_MAC_10_12);
	MAC_10_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_13, data_out=>output_MAC_10_13);
	MAC_10_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_14, data_out=>output_MAC_10_14);
	MAC_10_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_15, data_out=>output_MAC_10_15);
	MAC_10_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_16, data_out=>output_MAC_10_16);
	MAC_10_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_17, data_out=>output_MAC_10_17);
	MAC_10_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_18, data_out=>output_MAC_10_18);
	MAC_10_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_19, data_out=>output_MAC_10_19);
	MAC_10_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_20, data_out=>output_MAC_10_20);
	MAC_10_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_21, data_out=>output_MAC_10_21);
	MAC_10_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_22, data_out=>output_MAC_10_22);
	MAC_10_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_23, data_out=>output_MAC_10_23);
	MAC_10_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_24, data_out=>output_MAC_10_24);
	MAC_10_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_25, data_out=>output_MAC_10_25);
	MAC_10_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_26, data_out=>output_MAC_10_26);
	MAC_10_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_27, data_out=>output_MAC_10_27);
	MAC_10_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_28, data_out=>output_MAC_10_28);
	MAC_10_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_29, data_out=>output_MAC_10_29);
	MAC_10_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_30, data_out=>output_MAC_10_30);
	MAC_10_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_31, data_out=>output_MAC_10_31);
	MAC_11_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_0, data_out=>output_MAC_11_0);
	MAC_11_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_1, data_out=>output_MAC_11_1);
	MAC_11_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_2, data_out=>output_MAC_11_2);
	MAC_11_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_3, data_out=>output_MAC_11_3);
	MAC_11_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_4, data_out=>output_MAC_11_4);
	MAC_11_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_5, data_out=>output_MAC_11_5);
	MAC_11_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_6, data_out=>output_MAC_11_6);
	MAC_11_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_7, data_out=>output_MAC_11_7);
	MAC_11_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_8, data_out=>output_MAC_11_8);
	MAC_11_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_9, data_out=>output_MAC_11_9);
	MAC_11_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_10, data_out=>output_MAC_11_10);
	MAC_11_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_11, data_out=>output_MAC_11_11);
	MAC_11_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_12, data_out=>output_MAC_11_12);
	MAC_11_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_13, data_out=>output_MAC_11_13);
	MAC_11_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_14, data_out=>output_MAC_11_14);
	MAC_11_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_15, data_out=>output_MAC_11_15);
	MAC_11_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_16, data_out=>output_MAC_11_16);
	MAC_11_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_17, data_out=>output_MAC_11_17);
	MAC_11_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_18, data_out=>output_MAC_11_18);
	MAC_11_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_19, data_out=>output_MAC_11_19);
	MAC_11_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_20, data_out=>output_MAC_11_20);
	MAC_11_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_21, data_out=>output_MAC_11_21);
	MAC_11_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_22, data_out=>output_MAC_11_22);
	MAC_11_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_23, data_out=>output_MAC_11_23);
	MAC_11_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_24, data_out=>output_MAC_11_24);
	MAC_11_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_25, data_out=>output_MAC_11_25);
	MAC_11_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_26, data_out=>output_MAC_11_26);
	MAC_11_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_27, data_out=>output_MAC_11_27);
	MAC_11_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_28, data_out=>output_MAC_11_28);
	MAC_11_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_29, data_out=>output_MAC_11_29);
	MAC_11_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_30, data_out=>output_MAC_11_30);
	MAC_11_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_31, data_out=>output_MAC_11_31);
	MAC_12_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_0, data_out=>output_MAC_12_0);
	MAC_12_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_1, data_out=>output_MAC_12_1);
	MAC_12_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_2, data_out=>output_MAC_12_2);
	MAC_12_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_3, data_out=>output_MAC_12_3);
	MAC_12_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_4, data_out=>output_MAC_12_4);
	MAC_12_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_5, data_out=>output_MAC_12_5);
	MAC_12_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_6, data_out=>output_MAC_12_6);
	MAC_12_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_7, data_out=>output_MAC_12_7);
	MAC_12_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_8, data_out=>output_MAC_12_8);
	MAC_12_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_9, data_out=>output_MAC_12_9);
	MAC_12_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_10, data_out=>output_MAC_12_10);
	MAC_12_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_11, data_out=>output_MAC_12_11);
	MAC_12_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_12, data_out=>output_MAC_12_12);
	MAC_12_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_13, data_out=>output_MAC_12_13);
	MAC_12_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_14, data_out=>output_MAC_12_14);
	MAC_12_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_15, data_out=>output_MAC_12_15);
	MAC_12_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_16, data_out=>output_MAC_12_16);
	MAC_12_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_17, data_out=>output_MAC_12_17);
	MAC_12_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_18, data_out=>output_MAC_12_18);
	MAC_12_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_19, data_out=>output_MAC_12_19);
	MAC_12_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_20, data_out=>output_MAC_12_20);
	MAC_12_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_21, data_out=>output_MAC_12_21);
	MAC_12_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_22, data_out=>output_MAC_12_22);
	MAC_12_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_23, data_out=>output_MAC_12_23);
	MAC_12_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_24, data_out=>output_MAC_12_24);
	MAC_12_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_25, data_out=>output_MAC_12_25);
	MAC_12_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_26, data_out=>output_MAC_12_26);
	MAC_12_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_27, data_out=>output_MAC_12_27);
	MAC_12_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_28, data_out=>output_MAC_12_28);
	MAC_12_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_29, data_out=>output_MAC_12_29);
	MAC_12_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_30, data_out=>output_MAC_12_30);
	MAC_12_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_31, data_out=>output_MAC_12_31);
	MAC_13_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_0, data_out=>output_MAC_13_0);
	MAC_13_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_1, data_out=>output_MAC_13_1);
	MAC_13_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_2, data_out=>output_MAC_13_2);
	MAC_13_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_3, data_out=>output_MAC_13_3);
	MAC_13_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_4, data_out=>output_MAC_13_4);
	MAC_13_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_5, data_out=>output_MAC_13_5);
	MAC_13_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_6, data_out=>output_MAC_13_6);
	MAC_13_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_7, data_out=>output_MAC_13_7);
	MAC_13_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_8, data_out=>output_MAC_13_8);
	MAC_13_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_9, data_out=>output_MAC_13_9);
	MAC_13_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_10, data_out=>output_MAC_13_10);
	MAC_13_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_11, data_out=>output_MAC_13_11);
	MAC_13_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_12, data_out=>output_MAC_13_12);
	MAC_13_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_13, data_out=>output_MAC_13_13);
	MAC_13_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_14, data_out=>output_MAC_13_14);
	MAC_13_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_15, data_out=>output_MAC_13_15);
	MAC_13_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_16, data_out=>output_MAC_13_16);
	MAC_13_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_17, data_out=>output_MAC_13_17);
	MAC_13_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_18, data_out=>output_MAC_13_18);
	MAC_13_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_19, data_out=>output_MAC_13_19);
	MAC_13_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_20, data_out=>output_MAC_13_20);
	MAC_13_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_21, data_out=>output_MAC_13_21);
	MAC_13_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_22, data_out=>output_MAC_13_22);
	MAC_13_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_23, data_out=>output_MAC_13_23);
	MAC_13_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_24, data_out=>output_MAC_13_24);
	MAC_13_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_25, data_out=>output_MAC_13_25);
	MAC_13_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_26, data_out=>output_MAC_13_26);
	MAC_13_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_27, data_out=>output_MAC_13_27);
	MAC_13_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_28, data_out=>output_MAC_13_28);
	MAC_13_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_29, data_out=>output_MAC_13_29);
	MAC_13_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_30, data_out=>output_MAC_13_30);
	MAC_13_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_31, data_out=>output_MAC_13_31);
	MAC_14_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_0, data_out=>output_MAC_14_0);
	MAC_14_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_1, data_out=>output_MAC_14_1);
	MAC_14_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_2, data_out=>output_MAC_14_2);
	MAC_14_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_3, data_out=>output_MAC_14_3);
	MAC_14_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_4, data_out=>output_MAC_14_4);
	MAC_14_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_5, data_out=>output_MAC_14_5);
	MAC_14_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_6, data_out=>output_MAC_14_6);
	MAC_14_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_7, data_out=>output_MAC_14_7);
	MAC_14_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_8, data_out=>output_MAC_14_8);
	MAC_14_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_9, data_out=>output_MAC_14_9);
	MAC_14_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_10, data_out=>output_MAC_14_10);
	MAC_14_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_11, data_out=>output_MAC_14_11);
	MAC_14_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_12, data_out=>output_MAC_14_12);
	MAC_14_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_13, data_out=>output_MAC_14_13);
	MAC_14_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_14, data_out=>output_MAC_14_14);
	MAC_14_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_15, data_out=>output_MAC_14_15);
	MAC_14_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_16, data_out=>output_MAC_14_16);
	MAC_14_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_17, data_out=>output_MAC_14_17);
	MAC_14_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_18, data_out=>output_MAC_14_18);
	MAC_14_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_19, data_out=>output_MAC_14_19);
	MAC_14_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_20, data_out=>output_MAC_14_20);
	MAC_14_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_21, data_out=>output_MAC_14_21);
	MAC_14_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_22, data_out=>output_MAC_14_22);
	MAC_14_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_23, data_out=>output_MAC_14_23);
	MAC_14_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_24, data_out=>output_MAC_14_24);
	MAC_14_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_25, data_out=>output_MAC_14_25);
	MAC_14_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_26, data_out=>output_MAC_14_26);
	MAC_14_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_27, data_out=>output_MAC_14_27);
	MAC_14_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_28, data_out=>output_MAC_14_28);
	MAC_14_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_29, data_out=>output_MAC_14_29);
	MAC_14_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_30, data_out=>output_MAC_14_30);
	MAC_14_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_31, data_out=>output_MAC_14_31);
	MAC_15_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_0, data_out=>output_MAC_15_0);
	MAC_15_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_1, data_out=>output_MAC_15_1);
	MAC_15_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_2, data_out=>output_MAC_15_2);
	MAC_15_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_3, data_out=>output_MAC_15_3);
	MAC_15_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_4, data_out=>output_MAC_15_4);
	MAC_15_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_5, data_out=>output_MAC_15_5);
	MAC_15_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_6, data_out=>output_MAC_15_6);
	MAC_15_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_7, data_out=>output_MAC_15_7);
	MAC_15_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_8, data_out=>output_MAC_15_8);
	MAC_15_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_9, data_out=>output_MAC_15_9);
	MAC_15_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_10, data_out=>output_MAC_15_10);
	MAC_15_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_11, data_out=>output_MAC_15_11);
	MAC_15_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_12, data_out=>output_MAC_15_12);
	MAC_15_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_13, data_out=>output_MAC_15_13);
	MAC_15_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_14, data_out=>output_MAC_15_14);
	MAC_15_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_15, data_out=>output_MAC_15_15);
	MAC_15_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_16, data_out=>output_MAC_15_16);
	MAC_15_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_17, data_out=>output_MAC_15_17);
	MAC_15_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_18, data_out=>output_MAC_15_18);
	MAC_15_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_19, data_out=>output_MAC_15_19);
	MAC_15_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_20, data_out=>output_MAC_15_20);
	MAC_15_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_21, data_out=>output_MAC_15_21);
	MAC_15_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_22, data_out=>output_MAC_15_22);
	MAC_15_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_23, data_out=>output_MAC_15_23);
	MAC_15_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_24, data_out=>output_MAC_15_24);
	MAC_15_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_25, data_out=>output_MAC_15_25);
	MAC_15_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_26, data_out=>output_MAC_15_26);
	MAC_15_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_27, data_out=>output_MAC_15_27);
	MAC_15_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_28, data_out=>output_MAC_15_28);
	MAC_15_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_29, data_out=>output_MAC_15_29);
	MAC_15_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_30, data_out=>output_MAC_15_30);
	MAC_15_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_31, data_out=>output_MAC_15_31);
	MAC_16_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_0, data_out=>output_MAC_16_0);
	MAC_16_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_1, data_out=>output_MAC_16_1);
	MAC_16_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_2, data_out=>output_MAC_16_2);
	MAC_16_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_3, data_out=>output_MAC_16_3);
	MAC_16_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_4, data_out=>output_MAC_16_4);
	MAC_16_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_5, data_out=>output_MAC_16_5);
	MAC_16_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_6, data_out=>output_MAC_16_6);
	MAC_16_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_7, data_out=>output_MAC_16_7);
	MAC_16_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_8, data_out=>output_MAC_16_8);
	MAC_16_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_9, data_out=>output_MAC_16_9);
	MAC_16_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_10, data_out=>output_MAC_16_10);
	MAC_16_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_11, data_out=>output_MAC_16_11);
	MAC_16_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_12, data_out=>output_MAC_16_12);
	MAC_16_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_13, data_out=>output_MAC_16_13);
	MAC_16_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_14, data_out=>output_MAC_16_14);
	MAC_16_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_15, data_out=>output_MAC_16_15);
	MAC_16_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_16, data_out=>output_MAC_16_16);
	MAC_16_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_17, data_out=>output_MAC_16_17);
	MAC_16_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_18, data_out=>output_MAC_16_18);
	MAC_16_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_19, data_out=>output_MAC_16_19);
	MAC_16_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_20, data_out=>output_MAC_16_20);
	MAC_16_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_21, data_out=>output_MAC_16_21);
	MAC_16_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_22, data_out=>output_MAC_16_22);
	MAC_16_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_23, data_out=>output_MAC_16_23);
	MAC_16_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_24, data_out=>output_MAC_16_24);
	MAC_16_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_25, data_out=>output_MAC_16_25);
	MAC_16_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_26, data_out=>output_MAC_16_26);
	MAC_16_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_27, data_out=>output_MAC_16_27);
	MAC_16_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_28, data_out=>output_MAC_16_28);
	MAC_16_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_29, data_out=>output_MAC_16_29);
	MAC_16_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_30, data_out=>output_MAC_16_30);
	MAC_16_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_31, data_out=>output_MAC_16_31);
	MAC_17_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_0, data_out=>output_MAC_17_0);
	MAC_17_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_1, data_out=>output_MAC_17_1);
	MAC_17_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_2, data_out=>output_MAC_17_2);
	MAC_17_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_3, data_out=>output_MAC_17_3);
	MAC_17_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_4, data_out=>output_MAC_17_4);
	MAC_17_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_5, data_out=>output_MAC_17_5);
	MAC_17_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_6, data_out=>output_MAC_17_6);
	MAC_17_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_7, data_out=>output_MAC_17_7);
	MAC_17_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_8, data_out=>output_MAC_17_8);
	MAC_17_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_9, data_out=>output_MAC_17_9);
	MAC_17_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_10, data_out=>output_MAC_17_10);
	MAC_17_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_11, data_out=>output_MAC_17_11);
	MAC_17_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_12, data_out=>output_MAC_17_12);
	MAC_17_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_13, data_out=>output_MAC_17_13);
	MAC_17_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_14, data_out=>output_MAC_17_14);
	MAC_17_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_15, data_out=>output_MAC_17_15);
	MAC_17_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_16, data_out=>output_MAC_17_16);
	MAC_17_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_17, data_out=>output_MAC_17_17);
	MAC_17_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_18, data_out=>output_MAC_17_18);
	MAC_17_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_19, data_out=>output_MAC_17_19);
	MAC_17_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_20, data_out=>output_MAC_17_20);
	MAC_17_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_21, data_out=>output_MAC_17_21);
	MAC_17_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_22, data_out=>output_MAC_17_22);
	MAC_17_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_23, data_out=>output_MAC_17_23);
	MAC_17_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_24, data_out=>output_MAC_17_24);
	MAC_17_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_25, data_out=>output_MAC_17_25);
	MAC_17_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_26, data_out=>output_MAC_17_26);
	MAC_17_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_27, data_out=>output_MAC_17_27);
	MAC_17_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_28, data_out=>output_MAC_17_28);
	MAC_17_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_29, data_out=>output_MAC_17_29);
	MAC_17_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_30, data_out=>output_MAC_17_30);
	MAC_17_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_31, data_out=>output_MAC_17_31);
	MAC_18_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_0, data_out=>output_MAC_18_0);
	MAC_18_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_1, data_out=>output_MAC_18_1);
	MAC_18_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_2, data_out=>output_MAC_18_2);
	MAC_18_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_3, data_out=>output_MAC_18_3);
	MAC_18_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_4, data_out=>output_MAC_18_4);
	MAC_18_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_5, data_out=>output_MAC_18_5);
	MAC_18_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_6, data_out=>output_MAC_18_6);
	MAC_18_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_7, data_out=>output_MAC_18_7);
	MAC_18_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_8, data_out=>output_MAC_18_8);
	MAC_18_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_9, data_out=>output_MAC_18_9);
	MAC_18_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_10, data_out=>output_MAC_18_10);
	MAC_18_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_11, data_out=>output_MAC_18_11);
	MAC_18_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_12, data_out=>output_MAC_18_12);
	MAC_18_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_13, data_out=>output_MAC_18_13);
	MAC_18_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_14, data_out=>output_MAC_18_14);
	MAC_18_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_15, data_out=>output_MAC_18_15);
	MAC_18_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_16, data_out=>output_MAC_18_16);
	MAC_18_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_17, data_out=>output_MAC_18_17);
	MAC_18_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_18, data_out=>output_MAC_18_18);
	MAC_18_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_19, data_out=>output_MAC_18_19);
	MAC_18_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_20, data_out=>output_MAC_18_20);
	MAC_18_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_21, data_out=>output_MAC_18_21);
	MAC_18_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_22, data_out=>output_MAC_18_22);
	MAC_18_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_23, data_out=>output_MAC_18_23);
	MAC_18_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_24, data_out=>output_MAC_18_24);
	MAC_18_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_25, data_out=>output_MAC_18_25);
	MAC_18_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_26, data_out=>output_MAC_18_26);
	MAC_18_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_27, data_out=>output_MAC_18_27);
	MAC_18_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_28, data_out=>output_MAC_18_28);
	MAC_18_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_29, data_out=>output_MAC_18_29);
	MAC_18_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_30, data_out=>output_MAC_18_30);
	MAC_18_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_31, data_out=>output_MAC_18_31);
	MAC_19_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_0, data_out=>output_MAC_19_0);
	MAC_19_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_1, data_out=>output_MAC_19_1);
	MAC_19_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_2, data_out=>output_MAC_19_2);
	MAC_19_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_3, data_out=>output_MAC_19_3);
	MAC_19_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_4, data_out=>output_MAC_19_4);
	MAC_19_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_5, data_out=>output_MAC_19_5);
	MAC_19_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_6, data_out=>output_MAC_19_6);
	MAC_19_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_7, data_out=>output_MAC_19_7);
	MAC_19_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_8, data_out=>output_MAC_19_8);
	MAC_19_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_9, data_out=>output_MAC_19_9);
	MAC_19_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_10, data_out=>output_MAC_19_10);
	MAC_19_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_11, data_out=>output_MAC_19_11);
	MAC_19_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_12, data_out=>output_MAC_19_12);
	MAC_19_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_13, data_out=>output_MAC_19_13);
	MAC_19_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_14, data_out=>output_MAC_19_14);
	MAC_19_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_15, data_out=>output_MAC_19_15);
	MAC_19_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_16, data_out=>output_MAC_19_16);
	MAC_19_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_17, data_out=>output_MAC_19_17);
	MAC_19_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_18, data_out=>output_MAC_19_18);
	MAC_19_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_19, data_out=>output_MAC_19_19);
	MAC_19_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_20, data_out=>output_MAC_19_20);
	MAC_19_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_21, data_out=>output_MAC_19_21);
	MAC_19_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_22, data_out=>output_MAC_19_22);
	MAC_19_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_23, data_out=>output_MAC_19_23);
	MAC_19_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_24, data_out=>output_MAC_19_24);
	MAC_19_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_25, data_out=>output_MAC_19_25);
	MAC_19_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_26, data_out=>output_MAC_19_26);
	MAC_19_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_27, data_out=>output_MAC_19_27);
	MAC_19_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_28, data_out=>output_MAC_19_28);
	MAC_19_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_29, data_out=>output_MAC_19_29);
	MAC_19_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_30, data_out=>output_MAC_19_30);
	MAC_19_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_31, data_out=>output_MAC_19_31);
	MAC_20_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_0, data_out=>output_MAC_20_0);
	MAC_20_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_1, data_out=>output_MAC_20_1);
	MAC_20_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_2, data_out=>output_MAC_20_2);
	MAC_20_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_3, data_out=>output_MAC_20_3);
	MAC_20_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_4, data_out=>output_MAC_20_4);
	MAC_20_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_5, data_out=>output_MAC_20_5);
	MAC_20_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_6, data_out=>output_MAC_20_6);
	MAC_20_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_7, data_out=>output_MAC_20_7);
	MAC_20_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_8, data_out=>output_MAC_20_8);
	MAC_20_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_9, data_out=>output_MAC_20_9);
	MAC_20_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_10, data_out=>output_MAC_20_10);
	MAC_20_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_11, data_out=>output_MAC_20_11);
	MAC_20_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_12, data_out=>output_MAC_20_12);
	MAC_20_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_13, data_out=>output_MAC_20_13);
	MAC_20_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_14, data_out=>output_MAC_20_14);
	MAC_20_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_15, data_out=>output_MAC_20_15);
	MAC_20_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_16, data_out=>output_MAC_20_16);
	MAC_20_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_17, data_out=>output_MAC_20_17);
	MAC_20_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_18, data_out=>output_MAC_20_18);
	MAC_20_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_19, data_out=>output_MAC_20_19);
	MAC_20_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_20, data_out=>output_MAC_20_20);
	MAC_20_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_21, data_out=>output_MAC_20_21);
	MAC_20_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_22, data_out=>output_MAC_20_22);
	MAC_20_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_23, data_out=>output_MAC_20_23);
	MAC_20_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_24, data_out=>output_MAC_20_24);
	MAC_20_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_25, data_out=>output_MAC_20_25);
	MAC_20_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_26, data_out=>output_MAC_20_26);
	MAC_20_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_27, data_out=>output_MAC_20_27);
	MAC_20_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_28, data_out=>output_MAC_20_28);
	MAC_20_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_29, data_out=>output_MAC_20_29);
	MAC_20_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_30, data_out=>output_MAC_20_30);
	MAC_20_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_31, data_out=>output_MAC_20_31);
	MAC_21_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_0, data_out=>output_MAC_21_0);
	MAC_21_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_1, data_out=>output_MAC_21_1);
	MAC_21_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_2, data_out=>output_MAC_21_2);
	MAC_21_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_3, data_out=>output_MAC_21_3);
	MAC_21_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_4, data_out=>output_MAC_21_4);
	MAC_21_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_5, data_out=>output_MAC_21_5);
	MAC_21_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_6, data_out=>output_MAC_21_6);
	MAC_21_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_7, data_out=>output_MAC_21_7);
	MAC_21_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_8, data_out=>output_MAC_21_8);
	MAC_21_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_9, data_out=>output_MAC_21_9);
	MAC_21_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_10, data_out=>output_MAC_21_10);
	MAC_21_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_11, data_out=>output_MAC_21_11);
	MAC_21_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_12, data_out=>output_MAC_21_12);
	MAC_21_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_13, data_out=>output_MAC_21_13);
	MAC_21_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_14, data_out=>output_MAC_21_14);
	MAC_21_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_15, data_out=>output_MAC_21_15);
	MAC_21_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_16, data_out=>output_MAC_21_16);
	MAC_21_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_17, data_out=>output_MAC_21_17);
	MAC_21_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_18, data_out=>output_MAC_21_18);
	MAC_21_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_19, data_out=>output_MAC_21_19);
	MAC_21_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_20, data_out=>output_MAC_21_20);
	MAC_21_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_21, data_out=>output_MAC_21_21);
	MAC_21_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_22, data_out=>output_MAC_21_22);
	MAC_21_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_23, data_out=>output_MAC_21_23);
	MAC_21_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_24, data_out=>output_MAC_21_24);
	MAC_21_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_25, data_out=>output_MAC_21_25);
	MAC_21_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_26, data_out=>output_MAC_21_26);
	MAC_21_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_27, data_out=>output_MAC_21_27);
	MAC_21_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_28, data_out=>output_MAC_21_28);
	MAC_21_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_29, data_out=>output_MAC_21_29);
	MAC_21_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_30, data_out=>output_MAC_21_30);
	MAC_21_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_31, data_out=>output_MAC_21_31);
	MAC_22_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_0, data_out=>output_MAC_22_0);
	MAC_22_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_1, data_out=>output_MAC_22_1);
	MAC_22_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_2, data_out=>output_MAC_22_2);
	MAC_22_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_3, data_out=>output_MAC_22_3);
	MAC_22_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_4, data_out=>output_MAC_22_4);
	MAC_22_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_5, data_out=>output_MAC_22_5);
	MAC_22_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_6, data_out=>output_MAC_22_6);
	MAC_22_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_7, data_out=>output_MAC_22_7);
	MAC_22_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_8, data_out=>output_MAC_22_8);
	MAC_22_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_9, data_out=>output_MAC_22_9);
	MAC_22_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_10, data_out=>output_MAC_22_10);
	MAC_22_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_11, data_out=>output_MAC_22_11);
	MAC_22_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_12, data_out=>output_MAC_22_12);
	MAC_22_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_13, data_out=>output_MAC_22_13);
	MAC_22_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_14, data_out=>output_MAC_22_14);
	MAC_22_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_15, data_out=>output_MAC_22_15);
	MAC_22_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_16, data_out=>output_MAC_22_16);
	MAC_22_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_17, data_out=>output_MAC_22_17);
	MAC_22_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_18, data_out=>output_MAC_22_18);
	MAC_22_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_19, data_out=>output_MAC_22_19);
	MAC_22_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_20, data_out=>output_MAC_22_20);
	MAC_22_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_21, data_out=>output_MAC_22_21);
	MAC_22_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_22, data_out=>output_MAC_22_22);
	MAC_22_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_23, data_out=>output_MAC_22_23);
	MAC_22_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_24, data_out=>output_MAC_22_24);
	MAC_22_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_25, data_out=>output_MAC_22_25);
	MAC_22_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_26, data_out=>output_MAC_22_26);
	MAC_22_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_27, data_out=>output_MAC_22_27);
	MAC_22_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_28, data_out=>output_MAC_22_28);
	MAC_22_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_29, data_out=>output_MAC_22_29);
	MAC_22_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_30, data_out=>output_MAC_22_30);
	MAC_22_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_31, data_out=>output_MAC_22_31);
	MAC_23_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_0, data_out=>output_MAC_23_0);
	MAC_23_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_1, data_out=>output_MAC_23_1);
	MAC_23_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_2, data_out=>output_MAC_23_2);
	MAC_23_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_3, data_out=>output_MAC_23_3);
	MAC_23_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_4, data_out=>output_MAC_23_4);
	MAC_23_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_5, data_out=>output_MAC_23_5);
	MAC_23_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_6, data_out=>output_MAC_23_6);
	MAC_23_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_7, data_out=>output_MAC_23_7);
	MAC_23_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_8, data_out=>output_MAC_23_8);
	MAC_23_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_9, data_out=>output_MAC_23_9);
	MAC_23_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_10, data_out=>output_MAC_23_10);
	MAC_23_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_11, data_out=>output_MAC_23_11);
	MAC_23_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_12, data_out=>output_MAC_23_12);
	MAC_23_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_13, data_out=>output_MAC_23_13);
	MAC_23_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_14, data_out=>output_MAC_23_14);
	MAC_23_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_15, data_out=>output_MAC_23_15);
	MAC_23_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_16, data_out=>output_MAC_23_16);
	MAC_23_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_17, data_out=>output_MAC_23_17);
	MAC_23_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_18, data_out=>output_MAC_23_18);
	MAC_23_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_19, data_out=>output_MAC_23_19);
	MAC_23_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_20, data_out=>output_MAC_23_20);
	MAC_23_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_21, data_out=>output_MAC_23_21);
	MAC_23_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_22, data_out=>output_MAC_23_22);
	MAC_23_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_23, data_out=>output_MAC_23_23);
	MAC_23_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_24, data_out=>output_MAC_23_24);
	MAC_23_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_25, data_out=>output_MAC_23_25);
	MAC_23_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_26, data_out=>output_MAC_23_26);
	MAC_23_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_27, data_out=>output_MAC_23_27);
	MAC_23_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_28, data_out=>output_MAC_23_28);
	MAC_23_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_29, data_out=>output_MAC_23_29);
	MAC_23_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_30, data_out=>output_MAC_23_30);
	MAC_23_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_31, data_out=>output_MAC_23_31);
	MAC_24_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_0, data_out=>output_MAC_24_0);
	MAC_24_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_1, data_out=>output_MAC_24_1);
	MAC_24_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_2, data_out=>output_MAC_24_2);
	MAC_24_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_3, data_out=>output_MAC_24_3);
	MAC_24_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_4, data_out=>output_MAC_24_4);
	MAC_24_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_5, data_out=>output_MAC_24_5);
	MAC_24_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_6, data_out=>output_MAC_24_6);
	MAC_24_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_7, data_out=>output_MAC_24_7);
	MAC_24_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_8, data_out=>output_MAC_24_8);
	MAC_24_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_9, data_out=>output_MAC_24_9);
	MAC_24_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_10, data_out=>output_MAC_24_10);
	MAC_24_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_11, data_out=>output_MAC_24_11);
	MAC_24_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_12, data_out=>output_MAC_24_12);
	MAC_24_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_13, data_out=>output_MAC_24_13);
	MAC_24_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_14, data_out=>output_MAC_24_14);
	MAC_24_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_15, data_out=>output_MAC_24_15);
	MAC_24_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_16, data_out=>output_MAC_24_16);
	MAC_24_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_17, data_out=>output_MAC_24_17);
	MAC_24_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_18, data_out=>output_MAC_24_18);
	MAC_24_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_19, data_out=>output_MAC_24_19);
	MAC_24_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_20, data_out=>output_MAC_24_20);
	MAC_24_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_21, data_out=>output_MAC_24_21);
	MAC_24_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_22, data_out=>output_MAC_24_22);
	MAC_24_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_23, data_out=>output_MAC_24_23);
	MAC_24_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_24, data_out=>output_MAC_24_24);
	MAC_24_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_25, data_out=>output_MAC_24_25);
	MAC_24_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_26, data_out=>output_MAC_24_26);
	MAC_24_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_27, data_out=>output_MAC_24_27);
	MAC_24_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_28, data_out=>output_MAC_24_28);
	MAC_24_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_29, data_out=>output_MAC_24_29);
	MAC_24_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_30, data_out=>output_MAC_24_30);
	MAC_24_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_31, data_out=>output_MAC_24_31);
	MAC_25_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_0, data_out=>output_MAC_25_0);
	MAC_25_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_1, data_out=>output_MAC_25_1);
	MAC_25_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_2, data_out=>output_MAC_25_2);
	MAC_25_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_3, data_out=>output_MAC_25_3);
	MAC_25_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_4, data_out=>output_MAC_25_4);
	MAC_25_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_5, data_out=>output_MAC_25_5);
	MAC_25_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_6, data_out=>output_MAC_25_6);
	MAC_25_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_7, data_out=>output_MAC_25_7);
	MAC_25_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_8, data_out=>output_MAC_25_8);
	MAC_25_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_9, data_out=>output_MAC_25_9);
	MAC_25_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_10, data_out=>output_MAC_25_10);
	MAC_25_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_11, data_out=>output_MAC_25_11);
	MAC_25_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_12, data_out=>output_MAC_25_12);
	MAC_25_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_13, data_out=>output_MAC_25_13);
	MAC_25_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_14, data_out=>output_MAC_25_14);
	MAC_25_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_15, data_out=>output_MAC_25_15);
	MAC_25_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_16, data_out=>output_MAC_25_16);
	MAC_25_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_17, data_out=>output_MAC_25_17);
	MAC_25_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_18, data_out=>output_MAC_25_18);
	MAC_25_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_19, data_out=>output_MAC_25_19);
	MAC_25_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_20, data_out=>output_MAC_25_20);
	MAC_25_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_21, data_out=>output_MAC_25_21);
	MAC_25_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_22, data_out=>output_MAC_25_22);
	MAC_25_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_23, data_out=>output_MAC_25_23);
	MAC_25_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_24, data_out=>output_MAC_25_24);
	MAC_25_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_25, data_out=>output_MAC_25_25);
	MAC_25_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_26, data_out=>output_MAC_25_26);
	MAC_25_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_27, data_out=>output_MAC_25_27);
	MAC_25_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_28, data_out=>output_MAC_25_28);
	MAC_25_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_29, data_out=>output_MAC_25_29);
	MAC_25_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_30, data_out=>output_MAC_25_30);
	MAC_25_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_31, data_out=>output_MAC_25_31);
	MAC_26_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_0, data_out=>output_MAC_26_0);
	MAC_26_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_1, data_out=>output_MAC_26_1);
	MAC_26_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_2, data_out=>output_MAC_26_2);
	MAC_26_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_3, data_out=>output_MAC_26_3);
	MAC_26_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_4, data_out=>output_MAC_26_4);
	MAC_26_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_5, data_out=>output_MAC_26_5);
	MAC_26_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_6, data_out=>output_MAC_26_6);
	MAC_26_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_7, data_out=>output_MAC_26_7);
	MAC_26_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_8, data_out=>output_MAC_26_8);
	MAC_26_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_9, data_out=>output_MAC_26_9);
	MAC_26_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_10, data_out=>output_MAC_26_10);
	MAC_26_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_11, data_out=>output_MAC_26_11);
	MAC_26_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_12, data_out=>output_MAC_26_12);
	MAC_26_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_13, data_out=>output_MAC_26_13);
	MAC_26_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_14, data_out=>output_MAC_26_14);
	MAC_26_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_15, data_out=>output_MAC_26_15);
	MAC_26_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_16, data_out=>output_MAC_26_16);
	MAC_26_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_17, data_out=>output_MAC_26_17);
	MAC_26_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_18, data_out=>output_MAC_26_18);
	MAC_26_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_19, data_out=>output_MAC_26_19);
	MAC_26_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_20, data_out=>output_MAC_26_20);
	MAC_26_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_21, data_out=>output_MAC_26_21);
	MAC_26_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_22, data_out=>output_MAC_26_22);
	MAC_26_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_23, data_out=>output_MAC_26_23);
	MAC_26_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_24, data_out=>output_MAC_26_24);
	MAC_26_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_25, data_out=>output_MAC_26_25);
	MAC_26_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_26, data_out=>output_MAC_26_26);
	MAC_26_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_27, data_out=>output_MAC_26_27);
	MAC_26_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_28, data_out=>output_MAC_26_28);
	MAC_26_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_29, data_out=>output_MAC_26_29);
	MAC_26_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_30, data_out=>output_MAC_26_30);
	MAC_26_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_31, data_out=>output_MAC_26_31);
	MAC_27_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_0, data_out=>output_MAC_27_0);
	MAC_27_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_1, data_out=>output_MAC_27_1);
	MAC_27_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_2, data_out=>output_MAC_27_2);
	MAC_27_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_3, data_out=>output_MAC_27_3);
	MAC_27_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_4, data_out=>output_MAC_27_4);
	MAC_27_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_5, data_out=>output_MAC_27_5);
	MAC_27_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_6, data_out=>output_MAC_27_6);
	MAC_27_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_7, data_out=>output_MAC_27_7);
	MAC_27_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_8, data_out=>output_MAC_27_8);
	MAC_27_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_9, data_out=>output_MAC_27_9);
	MAC_27_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_10, data_out=>output_MAC_27_10);
	MAC_27_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_11, data_out=>output_MAC_27_11);
	MAC_27_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_12, data_out=>output_MAC_27_12);
	MAC_27_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_13, data_out=>output_MAC_27_13);
	MAC_27_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_14, data_out=>output_MAC_27_14);
	MAC_27_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_15, data_out=>output_MAC_27_15);
	MAC_27_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_16, data_out=>output_MAC_27_16);
	MAC_27_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_17, data_out=>output_MAC_27_17);
	MAC_27_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_18, data_out=>output_MAC_27_18);
	MAC_27_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_19, data_out=>output_MAC_27_19);
	MAC_27_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_20, data_out=>output_MAC_27_20);
	MAC_27_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_21, data_out=>output_MAC_27_21);
	MAC_27_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_22, data_out=>output_MAC_27_22);
	MAC_27_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_23, data_out=>output_MAC_27_23);
	MAC_27_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_24, data_out=>output_MAC_27_24);
	MAC_27_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_25, data_out=>output_MAC_27_25);
	MAC_27_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_26, data_out=>output_MAC_27_26);
	MAC_27_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_27, data_out=>output_MAC_27_27);
	MAC_27_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_28, data_out=>output_MAC_27_28);
	MAC_27_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_29, data_out=>output_MAC_27_29);
	MAC_27_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_30, data_out=>output_MAC_27_30);
	MAC_27_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_31, data_out=>output_MAC_27_31);
	MAC_28_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_0, data_out=>output_MAC_28_0);
	MAC_28_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_1, data_out=>output_MAC_28_1);
	MAC_28_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_2, data_out=>output_MAC_28_2);
	MAC_28_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_3, data_out=>output_MAC_28_3);
	MAC_28_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_4, data_out=>output_MAC_28_4);
	MAC_28_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_5, data_out=>output_MAC_28_5);
	MAC_28_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_6, data_out=>output_MAC_28_6);
	MAC_28_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_7, data_out=>output_MAC_28_7);
	MAC_28_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_8, data_out=>output_MAC_28_8);
	MAC_28_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_9, data_out=>output_MAC_28_9);
	MAC_28_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_10, data_out=>output_MAC_28_10);
	MAC_28_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_11, data_out=>output_MAC_28_11);
	MAC_28_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_12, data_out=>output_MAC_28_12);
	MAC_28_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_13, data_out=>output_MAC_28_13);
	MAC_28_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_14, data_out=>output_MAC_28_14);
	MAC_28_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_15, data_out=>output_MAC_28_15);
	MAC_28_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_16, data_out=>output_MAC_28_16);
	MAC_28_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_17, data_out=>output_MAC_28_17);
	MAC_28_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_18, data_out=>output_MAC_28_18);
	MAC_28_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_19, data_out=>output_MAC_28_19);
	MAC_28_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_20, data_out=>output_MAC_28_20);
	MAC_28_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_21, data_out=>output_MAC_28_21);
	MAC_28_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_22, data_out=>output_MAC_28_22);
	MAC_28_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_23, data_out=>output_MAC_28_23);
	MAC_28_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_24, data_out=>output_MAC_28_24);
	MAC_28_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_25, data_out=>output_MAC_28_25);
	MAC_28_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_26, data_out=>output_MAC_28_26);
	MAC_28_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_27, data_out=>output_MAC_28_27);
	MAC_28_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_28, data_out=>output_MAC_28_28);
	MAC_28_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_29, data_out=>output_MAC_28_29);
	MAC_28_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_30, data_out=>output_MAC_28_30);
	MAC_28_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_31, data_out=>output_MAC_28_31);
	MAC_29_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_0, data_out=>output_MAC_29_0);
	MAC_29_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_1, data_out=>output_MAC_29_1);
	MAC_29_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_2, data_out=>output_MAC_29_2);
	MAC_29_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_3, data_out=>output_MAC_29_3);
	MAC_29_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_4, data_out=>output_MAC_29_4);
	MAC_29_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_5, data_out=>output_MAC_29_5);
	MAC_29_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_6, data_out=>output_MAC_29_6);
	MAC_29_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_7, data_out=>output_MAC_29_7);
	MAC_29_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_8, data_out=>output_MAC_29_8);
	MAC_29_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_9, data_out=>output_MAC_29_9);
	MAC_29_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_10, data_out=>output_MAC_29_10);
	MAC_29_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_11, data_out=>output_MAC_29_11);
	MAC_29_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_12, data_out=>output_MAC_29_12);
	MAC_29_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_13, data_out=>output_MAC_29_13);
	MAC_29_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_14, data_out=>output_MAC_29_14);
	MAC_29_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_15, data_out=>output_MAC_29_15);
	MAC_29_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_16, data_out=>output_MAC_29_16);
	MAC_29_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_17, data_out=>output_MAC_29_17);
	MAC_29_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_18, data_out=>output_MAC_29_18);
	MAC_29_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_19, data_out=>output_MAC_29_19);
	MAC_29_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_20, data_out=>output_MAC_29_20);
	MAC_29_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_21, data_out=>output_MAC_29_21);
	MAC_29_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_22, data_out=>output_MAC_29_22);
	MAC_29_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_23, data_out=>output_MAC_29_23);
	MAC_29_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_24, data_out=>output_MAC_29_24);
	MAC_29_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_25, data_out=>output_MAC_29_25);
	MAC_29_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_26, data_out=>output_MAC_29_26);
	MAC_29_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_27, data_out=>output_MAC_29_27);
	MAC_29_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_28, data_out=>output_MAC_29_28);
	MAC_29_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_29, data_out=>output_MAC_29_29);
	MAC_29_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_30, data_out=>output_MAC_29_30);
	MAC_29_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_31, data_out=>output_MAC_29_31);
	MAC_30_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_0, data_out=>output_MAC_30_0);
	MAC_30_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_1, data_out=>output_MAC_30_1);
	MAC_30_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_2, data_out=>output_MAC_30_2);
	MAC_30_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_3, data_out=>output_MAC_30_3);
	MAC_30_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_4, data_out=>output_MAC_30_4);
	MAC_30_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_5, data_out=>output_MAC_30_5);
	MAC_30_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_6, data_out=>output_MAC_30_6);
	MAC_30_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_7, data_out=>output_MAC_30_7);
	MAC_30_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_8, data_out=>output_MAC_30_8);
	MAC_30_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_9, data_out=>output_MAC_30_9);
	MAC_30_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_10, data_out=>output_MAC_30_10);
	MAC_30_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_11, data_out=>output_MAC_30_11);
	MAC_30_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_12, data_out=>output_MAC_30_12);
	MAC_30_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_13, data_out=>output_MAC_30_13);
	MAC_30_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_14, data_out=>output_MAC_30_14);
	MAC_30_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_15, data_out=>output_MAC_30_15);
	MAC_30_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_16, data_out=>output_MAC_30_16);
	MAC_30_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_17, data_out=>output_MAC_30_17);
	MAC_30_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_18, data_out=>output_MAC_30_18);
	MAC_30_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_19, data_out=>output_MAC_30_19);
	MAC_30_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_20, data_out=>output_MAC_30_20);
	MAC_30_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_21, data_out=>output_MAC_30_21);
	MAC_30_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_22, data_out=>output_MAC_30_22);
	MAC_30_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_23, data_out=>output_MAC_30_23);
	MAC_30_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_24, data_out=>output_MAC_30_24);
	MAC_30_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_25, data_out=>output_MAC_30_25);
	MAC_30_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_26, data_out=>output_MAC_30_26);
	MAC_30_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_27, data_out=>output_MAC_30_27);
	MAC_30_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_28, data_out=>output_MAC_30_28);
	MAC_30_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_29, data_out=>output_MAC_30_29);
	MAC_30_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_30, data_out=>output_MAC_30_30);
	MAC_30_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_31, data_out=>output_MAC_30_31);
	MAC_31_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_0, data_out=>output_MAC_31_0);
	MAC_31_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_1, data_out=>output_MAC_31_1);
	MAC_31_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_2, data_out=>output_MAC_31_2);
	MAC_31_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_3, data_out=>output_MAC_31_3);
	MAC_31_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_4, data_out=>output_MAC_31_4);
	MAC_31_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_5, data_out=>output_MAC_31_5);
	MAC_31_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_6, data_out=>output_MAC_31_6);
	MAC_31_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_7, data_out=>output_MAC_31_7);
	MAC_31_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_8, data_out=>output_MAC_31_8);
	MAC_31_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_9, data_out=>output_MAC_31_9);
	MAC_31_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_10, data_out=>output_MAC_31_10);
	MAC_31_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_11, data_out=>output_MAC_31_11);
	MAC_31_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_12, data_out=>output_MAC_31_12);
	MAC_31_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_13, data_out=>output_MAC_31_13);
	MAC_31_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_14, data_out=>output_MAC_31_14);
	MAC_31_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_15, data_out=>output_MAC_31_15);
	MAC_31_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_16, data_out=>output_MAC_31_16);
	MAC_31_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_17, data_out=>output_MAC_31_17);
	MAC_31_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_18, data_out=>output_MAC_31_18);
	MAC_31_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_19, data_out=>output_MAC_31_19);
	MAC_31_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_20, data_out=>output_MAC_31_20);
	MAC_31_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_21, data_out=>output_MAC_31_21);
	MAC_31_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_22, data_out=>output_MAC_31_22);
	MAC_31_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_23, data_out=>output_MAC_31_23);
	MAC_31_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_24, data_out=>output_MAC_31_24);
	MAC_31_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_25, data_out=>output_MAC_31_25);
	MAC_31_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_26, data_out=>output_MAC_31_26);
	MAC_31_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_27, data_out=>output_MAC_31_27);
	MAC_31_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_28, data_out=>output_MAC_31_28);
	MAC_31_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_29, data_out=>output_MAC_31_29);
	MAC_31_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_30, data_out=>output_MAC_31_30);
	MAC_31_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_31, data_out=>output_MAC_31_31);
	MAC_32_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_0, data_out=>output_MAC_32_0);
	MAC_32_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_1, data_out=>output_MAC_32_1);
	MAC_32_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_2, data_out=>output_MAC_32_2);
	MAC_32_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_3, data_out=>output_MAC_32_3);
	MAC_32_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_4, data_out=>output_MAC_32_4);
	MAC_32_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_5, data_out=>output_MAC_32_5);
	MAC_32_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_6, data_out=>output_MAC_32_6);
	MAC_32_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_7, data_out=>output_MAC_32_7);
	MAC_32_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_8, data_out=>output_MAC_32_8);
	MAC_32_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_9, data_out=>output_MAC_32_9);
	MAC_32_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_10, data_out=>output_MAC_32_10);
	MAC_32_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_11, data_out=>output_MAC_32_11);
	MAC_32_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_12, data_out=>output_MAC_32_12);
	MAC_32_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_13, data_out=>output_MAC_32_13);
	MAC_32_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_14, data_out=>output_MAC_32_14);
	MAC_32_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_15, data_out=>output_MAC_32_15);
	MAC_32_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_16, data_out=>output_MAC_32_16);
	MAC_32_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_17, data_out=>output_MAC_32_17);
	MAC_32_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_18, data_out=>output_MAC_32_18);
	MAC_32_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_19, data_out=>output_MAC_32_19);
	MAC_32_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_20, data_out=>output_MAC_32_20);
	MAC_32_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_21, data_out=>output_MAC_32_21);
	MAC_32_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_22, data_out=>output_MAC_32_22);
	MAC_32_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_23, data_out=>output_MAC_32_23);
	MAC_32_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_24, data_out=>output_MAC_32_24);
	MAC_32_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_25, data_out=>output_MAC_32_25);
	MAC_32_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_26, data_out=>output_MAC_32_26);
	MAC_32_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_27, data_out=>output_MAC_32_27);
	MAC_32_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_28, data_out=>output_MAC_32_28);
	MAC_32_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_29, data_out=>output_MAC_32_29);
	MAC_32_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_30, data_out=>output_MAC_32_30);
	MAC_32_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_31, data_out=>output_MAC_32_31);
	MAC_33_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_0, data_out=>output_MAC_33_0);
	MAC_33_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_1, data_out=>output_MAC_33_1);
	MAC_33_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_2, data_out=>output_MAC_33_2);
	MAC_33_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_3, data_out=>output_MAC_33_3);
	MAC_33_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_4, data_out=>output_MAC_33_4);
	MAC_33_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_5, data_out=>output_MAC_33_5);
	MAC_33_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_6, data_out=>output_MAC_33_6);
	MAC_33_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_7, data_out=>output_MAC_33_7);
	MAC_33_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_8, data_out=>output_MAC_33_8);
	MAC_33_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_9, data_out=>output_MAC_33_9);
	MAC_33_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_10, data_out=>output_MAC_33_10);
	MAC_33_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_11, data_out=>output_MAC_33_11);
	MAC_33_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_12, data_out=>output_MAC_33_12);
	MAC_33_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_13, data_out=>output_MAC_33_13);
	MAC_33_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_14, data_out=>output_MAC_33_14);
	MAC_33_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_15, data_out=>output_MAC_33_15);
	MAC_33_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_16, data_out=>output_MAC_33_16);
	MAC_33_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_17, data_out=>output_MAC_33_17);
	MAC_33_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_18, data_out=>output_MAC_33_18);
	MAC_33_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_19, data_out=>output_MAC_33_19);
	MAC_33_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_20, data_out=>output_MAC_33_20);
	MAC_33_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_21, data_out=>output_MAC_33_21);
	MAC_33_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_22, data_out=>output_MAC_33_22);
	MAC_33_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_23, data_out=>output_MAC_33_23);
	MAC_33_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_24, data_out=>output_MAC_33_24);
	MAC_33_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_25, data_out=>output_MAC_33_25);
	MAC_33_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_26, data_out=>output_MAC_33_26);
	MAC_33_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_27, data_out=>output_MAC_33_27);
	MAC_33_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_28, data_out=>output_MAC_33_28);
	MAC_33_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_29, data_out=>output_MAC_33_29);
	MAC_33_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_30, data_out=>output_MAC_33_30);
	MAC_33_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_31, data_out=>output_MAC_33_31);
	MAC_34_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_0, data_out=>output_MAC_34_0);
	MAC_34_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_1, data_out=>output_MAC_34_1);
	MAC_34_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_2, data_out=>output_MAC_34_2);
	MAC_34_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_3, data_out=>output_MAC_34_3);
	MAC_34_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_4, data_out=>output_MAC_34_4);
	MAC_34_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_5, data_out=>output_MAC_34_5);
	MAC_34_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_6, data_out=>output_MAC_34_6);
	MAC_34_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_7, data_out=>output_MAC_34_7);
	MAC_34_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_8, data_out=>output_MAC_34_8);
	MAC_34_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_9, data_out=>output_MAC_34_9);
	MAC_34_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_10, data_out=>output_MAC_34_10);
	MAC_34_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_11, data_out=>output_MAC_34_11);
	MAC_34_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_12, data_out=>output_MAC_34_12);
	MAC_34_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_13, data_out=>output_MAC_34_13);
	MAC_34_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_14, data_out=>output_MAC_34_14);
	MAC_34_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_15, data_out=>output_MAC_34_15);
	MAC_34_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_16, data_out=>output_MAC_34_16);
	MAC_34_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_17, data_out=>output_MAC_34_17);
	MAC_34_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_18, data_out=>output_MAC_34_18);
	MAC_34_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_19, data_out=>output_MAC_34_19);
	MAC_34_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_20, data_out=>output_MAC_34_20);
	MAC_34_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_21, data_out=>output_MAC_34_21);
	MAC_34_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_22, data_out=>output_MAC_34_22);
	MAC_34_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_23, data_out=>output_MAC_34_23);
	MAC_34_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_24, data_out=>output_MAC_34_24);
	MAC_34_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_25, data_out=>output_MAC_34_25);
	MAC_34_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_26, data_out=>output_MAC_34_26);
	MAC_34_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_27, data_out=>output_MAC_34_27);
	MAC_34_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_28, data_out=>output_MAC_34_28);
	MAC_34_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_29, data_out=>output_MAC_34_29);
	MAC_34_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_30, data_out=>output_MAC_34_30);
	MAC_34_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_31, data_out=>output_MAC_34_31);
	MAC_35_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_0, data_out=>output_MAC_35_0);
	MAC_35_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_1, data_out=>output_MAC_35_1);
	MAC_35_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_2, data_out=>output_MAC_35_2);
	MAC_35_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_3, data_out=>output_MAC_35_3);
	MAC_35_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_4, data_out=>output_MAC_35_4);
	MAC_35_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_5, data_out=>output_MAC_35_5);
	MAC_35_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_6, data_out=>output_MAC_35_6);
	MAC_35_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_7, data_out=>output_MAC_35_7);
	MAC_35_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_8, data_out=>output_MAC_35_8);
	MAC_35_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_9, data_out=>output_MAC_35_9);
	MAC_35_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_10, data_out=>output_MAC_35_10);
	MAC_35_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_11, data_out=>output_MAC_35_11);
	MAC_35_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_12, data_out=>output_MAC_35_12);
	MAC_35_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_13, data_out=>output_MAC_35_13);
	MAC_35_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_14, data_out=>output_MAC_35_14);
	MAC_35_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_15, data_out=>output_MAC_35_15);
	MAC_35_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_16, data_out=>output_MAC_35_16);
	MAC_35_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_17, data_out=>output_MAC_35_17);
	MAC_35_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_18, data_out=>output_MAC_35_18);
	MAC_35_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_19, data_out=>output_MAC_35_19);
	MAC_35_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_20, data_out=>output_MAC_35_20);
	MAC_35_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_21, data_out=>output_MAC_35_21);
	MAC_35_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_22, data_out=>output_MAC_35_22);
	MAC_35_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_23, data_out=>output_MAC_35_23);
	MAC_35_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_24, data_out=>output_MAC_35_24);
	MAC_35_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_25, data_out=>output_MAC_35_25);
	MAC_35_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_26, data_out=>output_MAC_35_26);
	MAC_35_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_27, data_out=>output_MAC_35_27);
	MAC_35_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_28, data_out=>output_MAC_35_28);
	MAC_35_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_29, data_out=>output_MAC_35_29);
	MAC_35_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_30, data_out=>output_MAC_35_30);
	MAC_35_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_31, data_out=>output_MAC_35_31);
	MAC_36_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_0, data_out=>output_MAC_36_0);
	MAC_36_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_1, data_out=>output_MAC_36_1);
	MAC_36_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_2, data_out=>output_MAC_36_2);
	MAC_36_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_3, data_out=>output_MAC_36_3);
	MAC_36_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_4, data_out=>output_MAC_36_4);
	MAC_36_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_5, data_out=>output_MAC_36_5);
	MAC_36_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_6, data_out=>output_MAC_36_6);
	MAC_36_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_7, data_out=>output_MAC_36_7);
	MAC_36_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_8, data_out=>output_MAC_36_8);
	MAC_36_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_9, data_out=>output_MAC_36_9);
	MAC_36_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_10, data_out=>output_MAC_36_10);
	MAC_36_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_11, data_out=>output_MAC_36_11);
	MAC_36_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_12, data_out=>output_MAC_36_12);
	MAC_36_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_13, data_out=>output_MAC_36_13);
	MAC_36_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_14, data_out=>output_MAC_36_14);
	MAC_36_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_15, data_out=>output_MAC_36_15);
	MAC_36_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_16, data_out=>output_MAC_36_16);
	MAC_36_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_17, data_out=>output_MAC_36_17);
	MAC_36_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_18, data_out=>output_MAC_36_18);
	MAC_36_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_19, data_out=>output_MAC_36_19);
	MAC_36_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_20, data_out=>output_MAC_36_20);
	MAC_36_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_21, data_out=>output_MAC_36_21);
	MAC_36_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_22, data_out=>output_MAC_36_22);
	MAC_36_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_23, data_out=>output_MAC_36_23);
	MAC_36_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_24, data_out=>output_MAC_36_24);
	MAC_36_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_25, data_out=>output_MAC_36_25);
	MAC_36_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_26, data_out=>output_MAC_36_26);
	MAC_36_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_27, data_out=>output_MAC_36_27);
	MAC_36_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_28, data_out=>output_MAC_36_28);
	MAC_36_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_29, data_out=>output_MAC_36_29);
	MAC_36_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_30, data_out=>output_MAC_36_30);
	MAC_36_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_31, data_out=>output_MAC_36_31);
	MAC_37_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_0, data_out=>output_MAC_37_0);
	MAC_37_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_1, data_out=>output_MAC_37_1);
	MAC_37_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_2, data_out=>output_MAC_37_2);
	MAC_37_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_3, data_out=>output_MAC_37_3);
	MAC_37_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_4, data_out=>output_MAC_37_4);
	MAC_37_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_5, data_out=>output_MAC_37_5);
	MAC_37_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_6, data_out=>output_MAC_37_6);
	MAC_37_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_7, data_out=>output_MAC_37_7);
	MAC_37_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_8, data_out=>output_MAC_37_8);
	MAC_37_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_9, data_out=>output_MAC_37_9);
	MAC_37_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_10, data_out=>output_MAC_37_10);
	MAC_37_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_11, data_out=>output_MAC_37_11);
	MAC_37_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_12, data_out=>output_MAC_37_12);
	MAC_37_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_13, data_out=>output_MAC_37_13);
	MAC_37_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_14, data_out=>output_MAC_37_14);
	MAC_37_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_15, data_out=>output_MAC_37_15);
	MAC_37_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_16, data_out=>output_MAC_37_16);
	MAC_37_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_17, data_out=>output_MAC_37_17);
	MAC_37_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_18, data_out=>output_MAC_37_18);
	MAC_37_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_19, data_out=>output_MAC_37_19);
	MAC_37_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_20, data_out=>output_MAC_37_20);
	MAC_37_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_21, data_out=>output_MAC_37_21);
	MAC_37_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_22, data_out=>output_MAC_37_22);
	MAC_37_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_23, data_out=>output_MAC_37_23);
	MAC_37_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_24, data_out=>output_MAC_37_24);
	MAC_37_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_25, data_out=>output_MAC_37_25);
	MAC_37_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_26, data_out=>output_MAC_37_26);
	MAC_37_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_27, data_out=>output_MAC_37_27);
	MAC_37_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_28, data_out=>output_MAC_37_28);
	MAC_37_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_29, data_out=>output_MAC_37_29);
	MAC_37_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_30, data_out=>output_MAC_37_30);
	MAC_37_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_31, data_out=>output_MAC_37_31);
	MAC_38_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_0, data_out=>output_MAC_38_0);
	MAC_38_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_1, data_out=>output_MAC_38_1);
	MAC_38_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_2, data_out=>output_MAC_38_2);
	MAC_38_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_3, data_out=>output_MAC_38_3);
	MAC_38_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_4, data_out=>output_MAC_38_4);
	MAC_38_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_5, data_out=>output_MAC_38_5);
	MAC_38_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_6, data_out=>output_MAC_38_6);
	MAC_38_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_7, data_out=>output_MAC_38_7);
	MAC_38_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_8, data_out=>output_MAC_38_8);
	MAC_38_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_9, data_out=>output_MAC_38_9);
	MAC_38_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_10, data_out=>output_MAC_38_10);
	MAC_38_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_11, data_out=>output_MAC_38_11);
	MAC_38_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_12, data_out=>output_MAC_38_12);
	MAC_38_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_13, data_out=>output_MAC_38_13);
	MAC_38_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_14, data_out=>output_MAC_38_14);
	MAC_38_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_15, data_out=>output_MAC_38_15);
	MAC_38_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_16, data_out=>output_MAC_38_16);
	MAC_38_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_17, data_out=>output_MAC_38_17);
	MAC_38_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_18, data_out=>output_MAC_38_18);
	MAC_38_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_19, data_out=>output_MAC_38_19);
	MAC_38_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_20, data_out=>output_MAC_38_20);
	MAC_38_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_21, data_out=>output_MAC_38_21);
	MAC_38_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_22, data_out=>output_MAC_38_22);
	MAC_38_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_23, data_out=>output_MAC_38_23);
	MAC_38_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_24, data_out=>output_MAC_38_24);
	MAC_38_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_25, data_out=>output_MAC_38_25);
	MAC_38_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_26, data_out=>output_MAC_38_26);
	MAC_38_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_27, data_out=>output_MAC_38_27);
	MAC_38_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_28, data_out=>output_MAC_38_28);
	MAC_38_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_29, data_out=>output_MAC_38_29);
	MAC_38_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_30, data_out=>output_MAC_38_30);
	MAC_38_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_31, data_out=>output_MAC_38_31);
	MAC_39_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_0, data_out=>output_MAC_39_0);
	MAC_39_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_1, data_out=>output_MAC_39_1);
	MAC_39_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_2, data_out=>output_MAC_39_2);
	MAC_39_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_3, data_out=>output_MAC_39_3);
	MAC_39_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_4, data_out=>output_MAC_39_4);
	MAC_39_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_5, data_out=>output_MAC_39_5);
	MAC_39_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_6, data_out=>output_MAC_39_6);
	MAC_39_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_7, data_out=>output_MAC_39_7);
	MAC_39_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_8, data_out=>output_MAC_39_8);
	MAC_39_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_9, data_out=>output_MAC_39_9);
	MAC_39_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_10, data_out=>output_MAC_39_10);
	MAC_39_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_11, data_out=>output_MAC_39_11);
	MAC_39_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_12, data_out=>output_MAC_39_12);
	MAC_39_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_13, data_out=>output_MAC_39_13);
	MAC_39_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_14, data_out=>output_MAC_39_14);
	MAC_39_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_15, data_out=>output_MAC_39_15);
	MAC_39_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_16, data_out=>output_MAC_39_16);
	MAC_39_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_17, data_out=>output_MAC_39_17);
	MAC_39_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_18, data_out=>output_MAC_39_18);
	MAC_39_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_19, data_out=>output_MAC_39_19);
	MAC_39_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_20, data_out=>output_MAC_39_20);
	MAC_39_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_21, data_out=>output_MAC_39_21);
	MAC_39_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_22, data_out=>output_MAC_39_22);
	MAC_39_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_23, data_out=>output_MAC_39_23);
	MAC_39_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_24, data_out=>output_MAC_39_24);
	MAC_39_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_25, data_out=>output_MAC_39_25);
	MAC_39_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_26, data_out=>output_MAC_39_26);
	MAC_39_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_27, data_out=>output_MAC_39_27);
	MAC_39_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_28, data_out=>output_MAC_39_28);
	MAC_39_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_29, data_out=>output_MAC_39_29);
	MAC_39_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_30, data_out=>output_MAC_39_30);
	MAC_39_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_31, data_out=>output_MAC_39_31);
	MAC_40_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_0, data_out=>output_MAC_40_0);
	MAC_40_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_1, data_out=>output_MAC_40_1);
	MAC_40_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_2, data_out=>output_MAC_40_2);
	MAC_40_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_3, data_out=>output_MAC_40_3);
	MAC_40_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_4, data_out=>output_MAC_40_4);
	MAC_40_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_5, data_out=>output_MAC_40_5);
	MAC_40_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_6, data_out=>output_MAC_40_6);
	MAC_40_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_7, data_out=>output_MAC_40_7);
	MAC_40_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_8, data_out=>output_MAC_40_8);
	MAC_40_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_9, data_out=>output_MAC_40_9);
	MAC_40_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_10, data_out=>output_MAC_40_10);
	MAC_40_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_11, data_out=>output_MAC_40_11);
	MAC_40_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_12, data_out=>output_MAC_40_12);
	MAC_40_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_13, data_out=>output_MAC_40_13);
	MAC_40_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_14, data_out=>output_MAC_40_14);
	MAC_40_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_15, data_out=>output_MAC_40_15);
	MAC_40_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_16, data_out=>output_MAC_40_16);
	MAC_40_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_17, data_out=>output_MAC_40_17);
	MAC_40_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_18, data_out=>output_MAC_40_18);
	MAC_40_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_19, data_out=>output_MAC_40_19);
	MAC_40_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_20, data_out=>output_MAC_40_20);
	MAC_40_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_21, data_out=>output_MAC_40_21);
	MAC_40_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_22, data_out=>output_MAC_40_22);
	MAC_40_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_23, data_out=>output_MAC_40_23);
	MAC_40_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_24, data_out=>output_MAC_40_24);
	MAC_40_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_25, data_out=>output_MAC_40_25);
	MAC_40_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_26, data_out=>output_MAC_40_26);
	MAC_40_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_27, data_out=>output_MAC_40_27);
	MAC_40_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_28, data_out=>output_MAC_40_28);
	MAC_40_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_29, data_out=>output_MAC_40_29);
	MAC_40_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_30, data_out=>output_MAC_40_30);
	MAC_40_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_31, data_out=>output_MAC_40_31);
	MAC_41_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_0, data_out=>output_MAC_41_0);
	MAC_41_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_1, data_out=>output_MAC_41_1);
	MAC_41_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_2, data_out=>output_MAC_41_2);
	MAC_41_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_3, data_out=>output_MAC_41_3);
	MAC_41_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_4, data_out=>output_MAC_41_4);
	MAC_41_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_5, data_out=>output_MAC_41_5);
	MAC_41_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_6, data_out=>output_MAC_41_6);
	MAC_41_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_7, data_out=>output_MAC_41_7);
	MAC_41_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_8, data_out=>output_MAC_41_8);
	MAC_41_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_9, data_out=>output_MAC_41_9);
	MAC_41_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_10, data_out=>output_MAC_41_10);
	MAC_41_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_11, data_out=>output_MAC_41_11);
	MAC_41_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_12, data_out=>output_MAC_41_12);
	MAC_41_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_13, data_out=>output_MAC_41_13);
	MAC_41_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_14, data_out=>output_MAC_41_14);
	MAC_41_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_15, data_out=>output_MAC_41_15);
	MAC_41_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_16, data_out=>output_MAC_41_16);
	MAC_41_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_17, data_out=>output_MAC_41_17);
	MAC_41_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_18, data_out=>output_MAC_41_18);
	MAC_41_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_19, data_out=>output_MAC_41_19);
	MAC_41_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_20, data_out=>output_MAC_41_20);
	MAC_41_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_21, data_out=>output_MAC_41_21);
	MAC_41_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_22, data_out=>output_MAC_41_22);
	MAC_41_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_23, data_out=>output_MAC_41_23);
	MAC_41_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_24, data_out=>output_MAC_41_24);
	MAC_41_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_25, data_out=>output_MAC_41_25);
	MAC_41_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_26, data_out=>output_MAC_41_26);
	MAC_41_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_27, data_out=>output_MAC_41_27);
	MAC_41_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_28, data_out=>output_MAC_41_28);
	MAC_41_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_29, data_out=>output_MAC_41_29);
	MAC_41_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_30, data_out=>output_MAC_41_30);
	MAC_41_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_31, data_out=>output_MAC_41_31);
	MAC_42_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_0, data_out=>output_MAC_42_0);
	MAC_42_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_1, data_out=>output_MAC_42_1);
	MAC_42_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_2, data_out=>output_MAC_42_2);
	MAC_42_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_3, data_out=>output_MAC_42_3);
	MAC_42_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_4, data_out=>output_MAC_42_4);
	MAC_42_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_5, data_out=>output_MAC_42_5);
	MAC_42_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_6, data_out=>output_MAC_42_6);
	MAC_42_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_7, data_out=>output_MAC_42_7);
	MAC_42_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_8, data_out=>output_MAC_42_8);
	MAC_42_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_9, data_out=>output_MAC_42_9);
	MAC_42_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_10, data_out=>output_MAC_42_10);
	MAC_42_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_11, data_out=>output_MAC_42_11);
	MAC_42_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_12, data_out=>output_MAC_42_12);
	MAC_42_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_13, data_out=>output_MAC_42_13);
	MAC_42_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_14, data_out=>output_MAC_42_14);
	MAC_42_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_15, data_out=>output_MAC_42_15);
	MAC_42_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_16, data_out=>output_MAC_42_16);
	MAC_42_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_17, data_out=>output_MAC_42_17);
	MAC_42_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_18, data_out=>output_MAC_42_18);
	MAC_42_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_19, data_out=>output_MAC_42_19);
	MAC_42_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_20, data_out=>output_MAC_42_20);
	MAC_42_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_21, data_out=>output_MAC_42_21);
	MAC_42_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_22, data_out=>output_MAC_42_22);
	MAC_42_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_23, data_out=>output_MAC_42_23);
	MAC_42_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_24, data_out=>output_MAC_42_24);
	MAC_42_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_25, data_out=>output_MAC_42_25);
	MAC_42_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_26, data_out=>output_MAC_42_26);
	MAC_42_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_27, data_out=>output_MAC_42_27);
	MAC_42_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_28, data_out=>output_MAC_42_28);
	MAC_42_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_29, data_out=>output_MAC_42_29);
	MAC_42_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_30, data_out=>output_MAC_42_30);
	MAC_42_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_31, data_out=>output_MAC_42_31);
	MAC_43_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_0, data_out=>output_MAC_43_0);
	MAC_43_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_1, data_out=>output_MAC_43_1);
	MAC_43_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_2, data_out=>output_MAC_43_2);
	MAC_43_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_3, data_out=>output_MAC_43_3);
	MAC_43_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_4, data_out=>output_MAC_43_4);
	MAC_43_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_5, data_out=>output_MAC_43_5);
	MAC_43_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_6, data_out=>output_MAC_43_6);
	MAC_43_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_7, data_out=>output_MAC_43_7);
	MAC_43_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_8, data_out=>output_MAC_43_8);
	MAC_43_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_9, data_out=>output_MAC_43_9);
	MAC_43_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_10, data_out=>output_MAC_43_10);
	MAC_43_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_11, data_out=>output_MAC_43_11);
	MAC_43_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_12, data_out=>output_MAC_43_12);
	MAC_43_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_13, data_out=>output_MAC_43_13);
	MAC_43_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_14, data_out=>output_MAC_43_14);
	MAC_43_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_15, data_out=>output_MAC_43_15);
	MAC_43_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_16, data_out=>output_MAC_43_16);
	MAC_43_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_17, data_out=>output_MAC_43_17);
	MAC_43_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_18, data_out=>output_MAC_43_18);
	MAC_43_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_19, data_out=>output_MAC_43_19);
	MAC_43_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_20, data_out=>output_MAC_43_20);
	MAC_43_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_21, data_out=>output_MAC_43_21);
	MAC_43_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_22, data_out=>output_MAC_43_22);
	MAC_43_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_23, data_out=>output_MAC_43_23);
	MAC_43_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_24, data_out=>output_MAC_43_24);
	MAC_43_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_25, data_out=>output_MAC_43_25);
	MAC_43_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_26, data_out=>output_MAC_43_26);
	MAC_43_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_27, data_out=>output_MAC_43_27);
	MAC_43_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_28, data_out=>output_MAC_43_28);
	MAC_43_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_29, data_out=>output_MAC_43_29);
	MAC_43_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_30, data_out=>output_MAC_43_30);
	MAC_43_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_31, data_out=>output_MAC_43_31);
	MAC_44_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_0, data_out=>output_MAC_44_0);
	MAC_44_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_1, data_out=>output_MAC_44_1);
	MAC_44_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_2, data_out=>output_MAC_44_2);
	MAC_44_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_3, data_out=>output_MAC_44_3);
	MAC_44_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_4, data_out=>output_MAC_44_4);
	MAC_44_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_5, data_out=>output_MAC_44_5);
	MAC_44_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_6, data_out=>output_MAC_44_6);
	MAC_44_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_7, data_out=>output_MAC_44_7);
	MAC_44_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_8, data_out=>output_MAC_44_8);
	MAC_44_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_9, data_out=>output_MAC_44_9);
	MAC_44_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_10, data_out=>output_MAC_44_10);
	MAC_44_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_11, data_out=>output_MAC_44_11);
	MAC_44_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_12, data_out=>output_MAC_44_12);
	MAC_44_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_13, data_out=>output_MAC_44_13);
	MAC_44_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_14, data_out=>output_MAC_44_14);
	MAC_44_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_15, data_out=>output_MAC_44_15);
	MAC_44_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_16, data_out=>output_MAC_44_16);
	MAC_44_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_17, data_out=>output_MAC_44_17);
	MAC_44_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_18, data_out=>output_MAC_44_18);
	MAC_44_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_19, data_out=>output_MAC_44_19);
	MAC_44_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_20, data_out=>output_MAC_44_20);
	MAC_44_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_21, data_out=>output_MAC_44_21);
	MAC_44_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_22, data_out=>output_MAC_44_22);
	MAC_44_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_23, data_out=>output_MAC_44_23);
	MAC_44_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_24, data_out=>output_MAC_44_24);
	MAC_44_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_25, data_out=>output_MAC_44_25);
	MAC_44_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_26, data_out=>output_MAC_44_26);
	MAC_44_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_27, data_out=>output_MAC_44_27);
	MAC_44_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_28, data_out=>output_MAC_44_28);
	MAC_44_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_29, data_out=>output_MAC_44_29);
	MAC_44_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_30, data_out=>output_MAC_44_30);
	MAC_44_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_31, data_out=>output_MAC_44_31);
	MAC_45_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_0, data_out=>output_MAC_45_0);
	MAC_45_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_1, data_out=>output_MAC_45_1);
	MAC_45_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_2, data_out=>output_MAC_45_2);
	MAC_45_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_3, data_out=>output_MAC_45_3);
	MAC_45_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_4, data_out=>output_MAC_45_4);
	MAC_45_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_5, data_out=>output_MAC_45_5);
	MAC_45_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_6, data_out=>output_MAC_45_6);
	MAC_45_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_7, data_out=>output_MAC_45_7);
	MAC_45_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_8, data_out=>output_MAC_45_8);
	MAC_45_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_9, data_out=>output_MAC_45_9);
	MAC_45_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_10, data_out=>output_MAC_45_10);
	MAC_45_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_11, data_out=>output_MAC_45_11);
	MAC_45_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_12, data_out=>output_MAC_45_12);
	MAC_45_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_13, data_out=>output_MAC_45_13);
	MAC_45_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_14, data_out=>output_MAC_45_14);
	MAC_45_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_15, data_out=>output_MAC_45_15);
	MAC_45_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_16, data_out=>output_MAC_45_16);
	MAC_45_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_17, data_out=>output_MAC_45_17);
	MAC_45_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_18, data_out=>output_MAC_45_18);
	MAC_45_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_19, data_out=>output_MAC_45_19);
	MAC_45_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_20, data_out=>output_MAC_45_20);
	MAC_45_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_21, data_out=>output_MAC_45_21);
	MAC_45_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_22, data_out=>output_MAC_45_22);
	MAC_45_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_23, data_out=>output_MAC_45_23);
	MAC_45_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_24, data_out=>output_MAC_45_24);
	MAC_45_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_25, data_out=>output_MAC_45_25);
	MAC_45_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_26, data_out=>output_MAC_45_26);
	MAC_45_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_27, data_out=>output_MAC_45_27);
	MAC_45_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_28, data_out=>output_MAC_45_28);
	MAC_45_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_29, data_out=>output_MAC_45_29);
	MAC_45_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_30, data_out=>output_MAC_45_30);
	MAC_45_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_31, data_out=>output_MAC_45_31);
	MAC_46_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_0, data_out=>output_MAC_46_0);
	MAC_46_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_1, data_out=>output_MAC_46_1);
	MAC_46_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_2, data_out=>output_MAC_46_2);
	MAC_46_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_3, data_out=>output_MAC_46_3);
	MAC_46_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_4, data_out=>output_MAC_46_4);
	MAC_46_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_5, data_out=>output_MAC_46_5);
	MAC_46_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_6, data_out=>output_MAC_46_6);
	MAC_46_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_7, data_out=>output_MAC_46_7);
	MAC_46_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_8, data_out=>output_MAC_46_8);
	MAC_46_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_9, data_out=>output_MAC_46_9);
	MAC_46_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_10, data_out=>output_MAC_46_10);
	MAC_46_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_11, data_out=>output_MAC_46_11);
	MAC_46_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_12, data_out=>output_MAC_46_12);
	MAC_46_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_13, data_out=>output_MAC_46_13);
	MAC_46_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_14, data_out=>output_MAC_46_14);
	MAC_46_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_15, data_out=>output_MAC_46_15);
	MAC_46_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_16, data_out=>output_MAC_46_16);
	MAC_46_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_17, data_out=>output_MAC_46_17);
	MAC_46_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_18, data_out=>output_MAC_46_18);
	MAC_46_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_19, data_out=>output_MAC_46_19);
	MAC_46_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_20, data_out=>output_MAC_46_20);
	MAC_46_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_21, data_out=>output_MAC_46_21);
	MAC_46_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_22, data_out=>output_MAC_46_22);
	MAC_46_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_23, data_out=>output_MAC_46_23);
	MAC_46_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_24, data_out=>output_MAC_46_24);
	MAC_46_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_25, data_out=>output_MAC_46_25);
	MAC_46_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_26, data_out=>output_MAC_46_26);
	MAC_46_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_27, data_out=>output_MAC_46_27);
	MAC_46_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_28, data_out=>output_MAC_46_28);
	MAC_46_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_29, data_out=>output_MAC_46_29);
	MAC_46_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_30, data_out=>output_MAC_46_30);
	MAC_46_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_31, data_out=>output_MAC_46_31);
	MAC_47_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_0, data_out=>output_MAC_47_0);
	MAC_47_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_1, data_out=>output_MAC_47_1);
	MAC_47_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_2, data_out=>output_MAC_47_2);
	MAC_47_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_3, data_out=>output_MAC_47_3);
	MAC_47_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_4, data_out=>output_MAC_47_4);
	MAC_47_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_5, data_out=>output_MAC_47_5);
	MAC_47_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_6, data_out=>output_MAC_47_6);
	MAC_47_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_7, data_out=>output_MAC_47_7);
	MAC_47_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_8, data_out=>output_MAC_47_8);
	MAC_47_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_9, data_out=>output_MAC_47_9);
	MAC_47_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_10, data_out=>output_MAC_47_10);
	MAC_47_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_11, data_out=>output_MAC_47_11);
	MAC_47_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_12, data_out=>output_MAC_47_12);
	MAC_47_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_13, data_out=>output_MAC_47_13);
	MAC_47_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_14, data_out=>output_MAC_47_14);
	MAC_47_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_15, data_out=>output_MAC_47_15);
	MAC_47_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_16, data_out=>output_MAC_47_16);
	MAC_47_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_17, data_out=>output_MAC_47_17);
	MAC_47_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_18, data_out=>output_MAC_47_18);
	MAC_47_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_19, data_out=>output_MAC_47_19);
	MAC_47_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_20, data_out=>output_MAC_47_20);
	MAC_47_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_21, data_out=>output_MAC_47_21);
	MAC_47_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_22, data_out=>output_MAC_47_22);
	MAC_47_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_23, data_out=>output_MAC_47_23);
	MAC_47_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_24, data_out=>output_MAC_47_24);
	MAC_47_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_25, data_out=>output_MAC_47_25);
	MAC_47_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_26, data_out=>output_MAC_47_26);
	MAC_47_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_27, data_out=>output_MAC_47_27);
	MAC_47_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_28, data_out=>output_MAC_47_28);
	MAC_47_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_29, data_out=>output_MAC_47_29);
	MAC_47_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_30, data_out=>output_MAC_47_30);
	MAC_47_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_31, data_out=>output_MAC_47_31);
	MAC_48_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_0, data_out=>output_MAC_48_0);
	MAC_48_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_1, data_out=>output_MAC_48_1);
	MAC_48_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_2, data_out=>output_MAC_48_2);
	MAC_48_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_3, data_out=>output_MAC_48_3);
	MAC_48_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_4, data_out=>output_MAC_48_4);
	MAC_48_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_5, data_out=>output_MAC_48_5);
	MAC_48_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_6, data_out=>output_MAC_48_6);
	MAC_48_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_7, data_out=>output_MAC_48_7);
	MAC_48_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_8, data_out=>output_MAC_48_8);
	MAC_48_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_9, data_out=>output_MAC_48_9);
	MAC_48_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_10, data_out=>output_MAC_48_10);
	MAC_48_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_11, data_out=>output_MAC_48_11);
	MAC_48_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_12, data_out=>output_MAC_48_12);
	MAC_48_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_13, data_out=>output_MAC_48_13);
	MAC_48_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_14, data_out=>output_MAC_48_14);
	MAC_48_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_15, data_out=>output_MAC_48_15);
	MAC_48_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_16, data_out=>output_MAC_48_16);
	MAC_48_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_17, data_out=>output_MAC_48_17);
	MAC_48_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_18, data_out=>output_MAC_48_18);
	MAC_48_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_19, data_out=>output_MAC_48_19);
	MAC_48_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_20, data_out=>output_MAC_48_20);
	MAC_48_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_21, data_out=>output_MAC_48_21);
	MAC_48_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_22, data_out=>output_MAC_48_22);
	MAC_48_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_23, data_out=>output_MAC_48_23);
	MAC_48_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_24, data_out=>output_MAC_48_24);
	MAC_48_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_25, data_out=>output_MAC_48_25);
	MAC_48_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_26, data_out=>output_MAC_48_26);
	MAC_48_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_27, data_out=>output_MAC_48_27);
	MAC_48_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_28, data_out=>output_MAC_48_28);
	MAC_48_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_29, data_out=>output_MAC_48_29);
	MAC_48_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_30, data_out=>output_MAC_48_30);
	MAC_48_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_31, data_out=>output_MAC_48_31);
	MAC_49_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_0, data_out=>output_MAC_49_0);
	MAC_49_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_1, data_out=>output_MAC_49_1);
	MAC_49_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_2, data_out=>output_MAC_49_2);
	MAC_49_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_3, data_out=>output_MAC_49_3);
	MAC_49_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_4, data_out=>output_MAC_49_4);
	MAC_49_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_5, data_out=>output_MAC_49_5);
	MAC_49_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_6, data_out=>output_MAC_49_6);
	MAC_49_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_7, data_out=>output_MAC_49_7);
	MAC_49_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_8, data_out=>output_MAC_49_8);
	MAC_49_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_9, data_out=>output_MAC_49_9);
	MAC_49_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_10, data_out=>output_MAC_49_10);
	MAC_49_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_11, data_out=>output_MAC_49_11);
	MAC_49_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_12, data_out=>output_MAC_49_12);
	MAC_49_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_13, data_out=>output_MAC_49_13);
	MAC_49_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_14, data_out=>output_MAC_49_14);
	MAC_49_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_15, data_out=>output_MAC_49_15);
	MAC_49_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_16, data_out=>output_MAC_49_16);
	MAC_49_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_17, data_out=>output_MAC_49_17);
	MAC_49_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_18, data_out=>output_MAC_49_18);
	MAC_49_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_19, data_out=>output_MAC_49_19);
	MAC_49_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_20, data_out=>output_MAC_49_20);
	MAC_49_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_21, data_out=>output_MAC_49_21);
	MAC_49_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_22, data_out=>output_MAC_49_22);
	MAC_49_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_23, data_out=>output_MAC_49_23);
	MAC_49_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_24, data_out=>output_MAC_49_24);
	MAC_49_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_25, data_out=>output_MAC_49_25);
	MAC_49_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_26, data_out=>output_MAC_49_26);
	MAC_49_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_27, data_out=>output_MAC_49_27);
	MAC_49_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_28, data_out=>output_MAC_49_28);
	MAC_49_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_29, data_out=>output_MAC_49_29);
	MAC_49_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_30, data_out=>output_MAC_49_30);
	MAC_49_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_31, data_out=>output_MAC_49_31);
	MAC_50_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_0, data_out=>output_MAC_50_0);
	MAC_50_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_1, data_out=>output_MAC_50_1);
	MAC_50_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_2, data_out=>output_MAC_50_2);
	MAC_50_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_3, data_out=>output_MAC_50_3);
	MAC_50_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_4, data_out=>output_MAC_50_4);
	MAC_50_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_5, data_out=>output_MAC_50_5);
	MAC_50_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_6, data_out=>output_MAC_50_6);
	MAC_50_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_7, data_out=>output_MAC_50_7);
	MAC_50_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_8, data_out=>output_MAC_50_8);
	MAC_50_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_9, data_out=>output_MAC_50_9);
	MAC_50_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_10, data_out=>output_MAC_50_10);
	MAC_50_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_11, data_out=>output_MAC_50_11);
	MAC_50_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_12, data_out=>output_MAC_50_12);
	MAC_50_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_13, data_out=>output_MAC_50_13);
	MAC_50_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_14, data_out=>output_MAC_50_14);
	MAC_50_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_15, data_out=>output_MAC_50_15);
	MAC_50_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_16, data_out=>output_MAC_50_16);
	MAC_50_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_17, data_out=>output_MAC_50_17);
	MAC_50_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_18, data_out=>output_MAC_50_18);
	MAC_50_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_19, data_out=>output_MAC_50_19);
	MAC_50_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_20, data_out=>output_MAC_50_20);
	MAC_50_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_21, data_out=>output_MAC_50_21);
	MAC_50_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_22, data_out=>output_MAC_50_22);
	MAC_50_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_23, data_out=>output_MAC_50_23);
	MAC_50_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_24, data_out=>output_MAC_50_24);
	MAC_50_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_25, data_out=>output_MAC_50_25);
	MAC_50_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_26, data_out=>output_MAC_50_26);
	MAC_50_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_27, data_out=>output_MAC_50_27);
	MAC_50_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_28, data_out=>output_MAC_50_28);
	MAC_50_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_29, data_out=>output_MAC_50_29);
	MAC_50_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_30, data_out=>output_MAC_50_30);
	MAC_50_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_31, data_out=>output_MAC_50_31);
	MAC_51_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_0, data_out=>output_MAC_51_0);
	MAC_51_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_1, data_out=>output_MAC_51_1);
	MAC_51_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_2, data_out=>output_MAC_51_2);
	MAC_51_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_3, data_out=>output_MAC_51_3);
	MAC_51_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_4, data_out=>output_MAC_51_4);
	MAC_51_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_5, data_out=>output_MAC_51_5);
	MAC_51_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_6, data_out=>output_MAC_51_6);
	MAC_51_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_7, data_out=>output_MAC_51_7);
	MAC_51_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_8, data_out=>output_MAC_51_8);
	MAC_51_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_9, data_out=>output_MAC_51_9);
	MAC_51_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_10, data_out=>output_MAC_51_10);
	MAC_51_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_11, data_out=>output_MAC_51_11);
	MAC_51_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_12, data_out=>output_MAC_51_12);
	MAC_51_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_13, data_out=>output_MAC_51_13);
	MAC_51_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_14, data_out=>output_MAC_51_14);
	MAC_51_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_15, data_out=>output_MAC_51_15);
	MAC_51_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_16, data_out=>output_MAC_51_16);
	MAC_51_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_17, data_out=>output_MAC_51_17);
	MAC_51_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_18, data_out=>output_MAC_51_18);
	MAC_51_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_19, data_out=>output_MAC_51_19);
	MAC_51_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_20, data_out=>output_MAC_51_20);
	MAC_51_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_21, data_out=>output_MAC_51_21);
	MAC_51_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_22, data_out=>output_MAC_51_22);
	MAC_51_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_23, data_out=>output_MAC_51_23);
	MAC_51_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_24, data_out=>output_MAC_51_24);
	MAC_51_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_25, data_out=>output_MAC_51_25);
	MAC_51_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_26, data_out=>output_MAC_51_26);
	MAC_51_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_27, data_out=>output_MAC_51_27);
	MAC_51_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_28, data_out=>output_MAC_51_28);
	MAC_51_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_29, data_out=>output_MAC_51_29);
	MAC_51_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_30, data_out=>output_MAC_51_30);
	MAC_51_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_31, data_out=>output_MAC_51_31);
	MAC_52_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_0, data_out=>output_MAC_52_0);
	MAC_52_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_1, data_out=>output_MAC_52_1);
	MAC_52_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_2, data_out=>output_MAC_52_2);
	MAC_52_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_3, data_out=>output_MAC_52_3);
	MAC_52_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_4, data_out=>output_MAC_52_4);
	MAC_52_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_5, data_out=>output_MAC_52_5);
	MAC_52_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_6, data_out=>output_MAC_52_6);
	MAC_52_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_7, data_out=>output_MAC_52_7);
	MAC_52_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_8, data_out=>output_MAC_52_8);
	MAC_52_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_9, data_out=>output_MAC_52_9);
	MAC_52_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_10, data_out=>output_MAC_52_10);
	MAC_52_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_11, data_out=>output_MAC_52_11);
	MAC_52_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_12, data_out=>output_MAC_52_12);
	MAC_52_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_13, data_out=>output_MAC_52_13);
	MAC_52_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_14, data_out=>output_MAC_52_14);
	MAC_52_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_15, data_out=>output_MAC_52_15);
	MAC_52_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_16, data_out=>output_MAC_52_16);
	MAC_52_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_17, data_out=>output_MAC_52_17);
	MAC_52_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_18, data_out=>output_MAC_52_18);
	MAC_52_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_19, data_out=>output_MAC_52_19);
	MAC_52_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_20, data_out=>output_MAC_52_20);
	MAC_52_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_21, data_out=>output_MAC_52_21);
	MAC_52_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_22, data_out=>output_MAC_52_22);
	MAC_52_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_23, data_out=>output_MAC_52_23);
	MAC_52_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_24, data_out=>output_MAC_52_24);
	MAC_52_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_25, data_out=>output_MAC_52_25);
	MAC_52_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_26, data_out=>output_MAC_52_26);
	MAC_52_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_27, data_out=>output_MAC_52_27);
	MAC_52_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_28, data_out=>output_MAC_52_28);
	MAC_52_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_29, data_out=>output_MAC_52_29);
	MAC_52_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_30, data_out=>output_MAC_52_30);
	MAC_52_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_31, data_out=>output_MAC_52_31);
	MAC_53_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_0, data_out=>output_MAC_53_0);
	MAC_53_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_1, data_out=>output_MAC_53_1);
	MAC_53_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_2, data_out=>output_MAC_53_2);
	MAC_53_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_3, data_out=>output_MAC_53_3);
	MAC_53_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_4, data_out=>output_MAC_53_4);
	MAC_53_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_5, data_out=>output_MAC_53_5);
	MAC_53_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_6, data_out=>output_MAC_53_6);
	MAC_53_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_7, data_out=>output_MAC_53_7);
	MAC_53_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_8, data_out=>output_MAC_53_8);
	MAC_53_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_9, data_out=>output_MAC_53_9);
	MAC_53_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_10, data_out=>output_MAC_53_10);
	MAC_53_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_11, data_out=>output_MAC_53_11);
	MAC_53_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_12, data_out=>output_MAC_53_12);
	MAC_53_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_13, data_out=>output_MAC_53_13);
	MAC_53_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_14, data_out=>output_MAC_53_14);
	MAC_53_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_15, data_out=>output_MAC_53_15);
	MAC_53_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_16, data_out=>output_MAC_53_16);
	MAC_53_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_17, data_out=>output_MAC_53_17);
	MAC_53_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_18, data_out=>output_MAC_53_18);
	MAC_53_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_19, data_out=>output_MAC_53_19);
	MAC_53_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_20, data_out=>output_MAC_53_20);
	MAC_53_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_21, data_out=>output_MAC_53_21);
	MAC_53_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_22, data_out=>output_MAC_53_22);
	MAC_53_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_23, data_out=>output_MAC_53_23);
	MAC_53_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_24, data_out=>output_MAC_53_24);
	MAC_53_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_25, data_out=>output_MAC_53_25);
	MAC_53_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_26, data_out=>output_MAC_53_26);
	MAC_53_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_27, data_out=>output_MAC_53_27);
	MAC_53_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_28, data_out=>output_MAC_53_28);
	MAC_53_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_29, data_out=>output_MAC_53_29);
	MAC_53_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_30, data_out=>output_MAC_53_30);
	MAC_53_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_31, data_out=>output_MAC_53_31);
	MAC_54_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_0, data_out=>output_MAC_54_0);
	MAC_54_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_1, data_out=>output_MAC_54_1);
	MAC_54_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_2, data_out=>output_MAC_54_2);
	MAC_54_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_3, data_out=>output_MAC_54_3);
	MAC_54_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_4, data_out=>output_MAC_54_4);
	MAC_54_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_5, data_out=>output_MAC_54_5);
	MAC_54_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_6, data_out=>output_MAC_54_6);
	MAC_54_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_7, data_out=>output_MAC_54_7);
	MAC_54_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_8, data_out=>output_MAC_54_8);
	MAC_54_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_9, data_out=>output_MAC_54_9);
	MAC_54_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_10, data_out=>output_MAC_54_10);
	MAC_54_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_11, data_out=>output_MAC_54_11);
	MAC_54_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_12, data_out=>output_MAC_54_12);
	MAC_54_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_13, data_out=>output_MAC_54_13);
	MAC_54_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_14, data_out=>output_MAC_54_14);
	MAC_54_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_15, data_out=>output_MAC_54_15);
	MAC_54_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_16, data_out=>output_MAC_54_16);
	MAC_54_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_17, data_out=>output_MAC_54_17);
	MAC_54_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_18, data_out=>output_MAC_54_18);
	MAC_54_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_19, data_out=>output_MAC_54_19);
	MAC_54_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_20, data_out=>output_MAC_54_20);
	MAC_54_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_21, data_out=>output_MAC_54_21);
	MAC_54_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_22, data_out=>output_MAC_54_22);
	MAC_54_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_23, data_out=>output_MAC_54_23);
	MAC_54_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_24, data_out=>output_MAC_54_24);
	MAC_54_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_25, data_out=>output_MAC_54_25);
	MAC_54_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_26, data_out=>output_MAC_54_26);
	MAC_54_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_27, data_out=>output_MAC_54_27);
	MAC_54_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_28, data_out=>output_MAC_54_28);
	MAC_54_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_29, data_out=>output_MAC_54_29);
	MAC_54_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_30, data_out=>output_MAC_54_30);
	MAC_54_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_31, data_out=>output_MAC_54_31);
	MAC_55_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_0, data_out=>output_MAC_55_0);
	MAC_55_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_1, data_out=>output_MAC_55_1);
	MAC_55_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_2, data_out=>output_MAC_55_2);
	MAC_55_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_3, data_out=>output_MAC_55_3);
	MAC_55_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_4, data_out=>output_MAC_55_4);
	MAC_55_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_5, data_out=>output_MAC_55_5);
	MAC_55_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_6, data_out=>output_MAC_55_6);
	MAC_55_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_7, data_out=>output_MAC_55_7);
	MAC_55_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_8, data_out=>output_MAC_55_8);
	MAC_55_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_9, data_out=>output_MAC_55_9);
	MAC_55_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_10, data_out=>output_MAC_55_10);
	MAC_55_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_11, data_out=>output_MAC_55_11);
	MAC_55_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_12, data_out=>output_MAC_55_12);
	MAC_55_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_13, data_out=>output_MAC_55_13);
	MAC_55_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_14, data_out=>output_MAC_55_14);
	MAC_55_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_15, data_out=>output_MAC_55_15);
	MAC_55_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_16, data_out=>output_MAC_55_16);
	MAC_55_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_17, data_out=>output_MAC_55_17);
	MAC_55_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_18, data_out=>output_MAC_55_18);
	MAC_55_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_19, data_out=>output_MAC_55_19);
	MAC_55_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_20, data_out=>output_MAC_55_20);
	MAC_55_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_21, data_out=>output_MAC_55_21);
	MAC_55_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_22, data_out=>output_MAC_55_22);
	MAC_55_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_23, data_out=>output_MAC_55_23);
	MAC_55_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_24, data_out=>output_MAC_55_24);
	MAC_55_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_25, data_out=>output_MAC_55_25);
	MAC_55_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_26, data_out=>output_MAC_55_26);
	MAC_55_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_27, data_out=>output_MAC_55_27);
	MAC_55_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_28, data_out=>output_MAC_55_28);
	MAC_55_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_29, data_out=>output_MAC_55_29);
	MAC_55_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_30, data_out=>output_MAC_55_30);
	MAC_55_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_31, data_out=>output_MAC_55_31);
	MAC_56_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_0, data_out=>output_MAC_56_0);
	MAC_56_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_1, data_out=>output_MAC_56_1);
	MAC_56_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_2, data_out=>output_MAC_56_2);
	MAC_56_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_3, data_out=>output_MAC_56_3);
	MAC_56_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_4, data_out=>output_MAC_56_4);
	MAC_56_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_5, data_out=>output_MAC_56_5);
	MAC_56_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_6, data_out=>output_MAC_56_6);
	MAC_56_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_7, data_out=>output_MAC_56_7);
	MAC_56_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_8, data_out=>output_MAC_56_8);
	MAC_56_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_9, data_out=>output_MAC_56_9);
	MAC_56_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_10, data_out=>output_MAC_56_10);
	MAC_56_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_11, data_out=>output_MAC_56_11);
	MAC_56_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_12, data_out=>output_MAC_56_12);
	MAC_56_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_13, data_out=>output_MAC_56_13);
	MAC_56_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_14, data_out=>output_MAC_56_14);
	MAC_56_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_15, data_out=>output_MAC_56_15);
	MAC_56_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_16, data_out=>output_MAC_56_16);
	MAC_56_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_17, data_out=>output_MAC_56_17);
	MAC_56_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_18, data_out=>output_MAC_56_18);
	MAC_56_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_19, data_out=>output_MAC_56_19);
	MAC_56_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_20, data_out=>output_MAC_56_20);
	MAC_56_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_21, data_out=>output_MAC_56_21);
	MAC_56_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_22, data_out=>output_MAC_56_22);
	MAC_56_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_23, data_out=>output_MAC_56_23);
	MAC_56_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_24, data_out=>output_MAC_56_24);
	MAC_56_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_25, data_out=>output_MAC_56_25);
	MAC_56_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_26, data_out=>output_MAC_56_26);
	MAC_56_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_27, data_out=>output_MAC_56_27);
	MAC_56_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_28, data_out=>output_MAC_56_28);
	MAC_56_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_29, data_out=>output_MAC_56_29);
	MAC_56_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_30, data_out=>output_MAC_56_30);
	MAC_56_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_31, data_out=>output_MAC_56_31);
	MAC_57_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_0, data_out=>output_MAC_57_0);
	MAC_57_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_1, data_out=>output_MAC_57_1);
	MAC_57_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_2, data_out=>output_MAC_57_2);
	MAC_57_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_3, data_out=>output_MAC_57_3);
	MAC_57_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_4, data_out=>output_MAC_57_4);
	MAC_57_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_5, data_out=>output_MAC_57_5);
	MAC_57_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_6, data_out=>output_MAC_57_6);
	MAC_57_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_7, data_out=>output_MAC_57_7);
	MAC_57_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_8, data_out=>output_MAC_57_8);
	MAC_57_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_9, data_out=>output_MAC_57_9);
	MAC_57_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_10, data_out=>output_MAC_57_10);
	MAC_57_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_11, data_out=>output_MAC_57_11);
	MAC_57_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_12, data_out=>output_MAC_57_12);
	MAC_57_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_13, data_out=>output_MAC_57_13);
	MAC_57_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_14, data_out=>output_MAC_57_14);
	MAC_57_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_15, data_out=>output_MAC_57_15);
	MAC_57_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_16, data_out=>output_MAC_57_16);
	MAC_57_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_17, data_out=>output_MAC_57_17);
	MAC_57_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_18, data_out=>output_MAC_57_18);
	MAC_57_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_19, data_out=>output_MAC_57_19);
	MAC_57_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_20, data_out=>output_MAC_57_20);
	MAC_57_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_21, data_out=>output_MAC_57_21);
	MAC_57_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_22, data_out=>output_MAC_57_22);
	MAC_57_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_23, data_out=>output_MAC_57_23);
	MAC_57_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_24, data_out=>output_MAC_57_24);
	MAC_57_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_25, data_out=>output_MAC_57_25);
	MAC_57_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_26, data_out=>output_MAC_57_26);
	MAC_57_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_27, data_out=>output_MAC_57_27);
	MAC_57_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_28, data_out=>output_MAC_57_28);
	MAC_57_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_29, data_out=>output_MAC_57_29);
	MAC_57_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_30, data_out=>output_MAC_57_30);
	MAC_57_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_31, data_out=>output_MAC_57_31);
	MAC_58_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_0, data_out=>output_MAC_58_0);
	MAC_58_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_1, data_out=>output_MAC_58_1);
	MAC_58_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_2, data_out=>output_MAC_58_2);
	MAC_58_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_3, data_out=>output_MAC_58_3);
	MAC_58_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_4, data_out=>output_MAC_58_4);
	MAC_58_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_5, data_out=>output_MAC_58_5);
	MAC_58_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_6, data_out=>output_MAC_58_6);
	MAC_58_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_7, data_out=>output_MAC_58_7);
	MAC_58_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_8, data_out=>output_MAC_58_8);
	MAC_58_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_9, data_out=>output_MAC_58_9);
	MAC_58_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_10, data_out=>output_MAC_58_10);
	MAC_58_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_11, data_out=>output_MAC_58_11);
	MAC_58_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_12, data_out=>output_MAC_58_12);
	MAC_58_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_13, data_out=>output_MAC_58_13);
	MAC_58_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_14, data_out=>output_MAC_58_14);
	MAC_58_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_15, data_out=>output_MAC_58_15);
	MAC_58_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_16, data_out=>output_MAC_58_16);
	MAC_58_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_17, data_out=>output_MAC_58_17);
	MAC_58_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_18, data_out=>output_MAC_58_18);
	MAC_58_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_19, data_out=>output_MAC_58_19);
	MAC_58_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_20, data_out=>output_MAC_58_20);
	MAC_58_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_21, data_out=>output_MAC_58_21);
	MAC_58_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_22, data_out=>output_MAC_58_22);
	MAC_58_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_23, data_out=>output_MAC_58_23);
	MAC_58_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_24, data_out=>output_MAC_58_24);
	MAC_58_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_25, data_out=>output_MAC_58_25);
	MAC_58_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_26, data_out=>output_MAC_58_26);
	MAC_58_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_27, data_out=>output_MAC_58_27);
	MAC_58_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_28, data_out=>output_MAC_58_28);
	MAC_58_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_29, data_out=>output_MAC_58_29);
	MAC_58_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_30, data_out=>output_MAC_58_30);
	MAC_58_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_31, data_out=>output_MAC_58_31);
	MAC_59_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_0, data_out=>output_MAC_59_0);
	MAC_59_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_1, data_out=>output_MAC_59_1);
	MAC_59_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_2, data_out=>output_MAC_59_2);
	MAC_59_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_3, data_out=>output_MAC_59_3);
	MAC_59_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_4, data_out=>output_MAC_59_4);
	MAC_59_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_5, data_out=>output_MAC_59_5);
	MAC_59_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_6, data_out=>output_MAC_59_6);
	MAC_59_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_7, data_out=>output_MAC_59_7);
	MAC_59_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_8, data_out=>output_MAC_59_8);
	MAC_59_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_9, data_out=>output_MAC_59_9);
	MAC_59_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_10, data_out=>output_MAC_59_10);
	MAC_59_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_11, data_out=>output_MAC_59_11);
	MAC_59_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_12, data_out=>output_MAC_59_12);
	MAC_59_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_13, data_out=>output_MAC_59_13);
	MAC_59_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_14, data_out=>output_MAC_59_14);
	MAC_59_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_15, data_out=>output_MAC_59_15);
	MAC_59_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_16, data_out=>output_MAC_59_16);
	MAC_59_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_17, data_out=>output_MAC_59_17);
	MAC_59_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_18, data_out=>output_MAC_59_18);
	MAC_59_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_19, data_out=>output_MAC_59_19);
	MAC_59_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_20, data_out=>output_MAC_59_20);
	MAC_59_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_21, data_out=>output_MAC_59_21);
	MAC_59_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_22, data_out=>output_MAC_59_22);
	MAC_59_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_23, data_out=>output_MAC_59_23);
	MAC_59_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_24, data_out=>output_MAC_59_24);
	MAC_59_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_25, data_out=>output_MAC_59_25);
	MAC_59_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_26, data_out=>output_MAC_59_26);
	MAC_59_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_27, data_out=>output_MAC_59_27);
	MAC_59_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_28, data_out=>output_MAC_59_28);
	MAC_59_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_29, data_out=>output_MAC_59_29);
	MAC_59_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_30, data_out=>output_MAC_59_30);
	MAC_59_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_31, data_out=>output_MAC_59_31);
	MAC_60_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_0, data_out=>output_MAC_60_0);
	MAC_60_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_1, data_out=>output_MAC_60_1);
	MAC_60_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_2, data_out=>output_MAC_60_2);
	MAC_60_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_3, data_out=>output_MAC_60_3);
	MAC_60_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_4, data_out=>output_MAC_60_4);
	MAC_60_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_5, data_out=>output_MAC_60_5);
	MAC_60_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_6, data_out=>output_MAC_60_6);
	MAC_60_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_7, data_out=>output_MAC_60_7);
	MAC_60_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_8, data_out=>output_MAC_60_8);
	MAC_60_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_9, data_out=>output_MAC_60_9);
	MAC_60_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_10, data_out=>output_MAC_60_10);
	MAC_60_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_11, data_out=>output_MAC_60_11);
	MAC_60_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_12, data_out=>output_MAC_60_12);
	MAC_60_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_13, data_out=>output_MAC_60_13);
	MAC_60_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_14, data_out=>output_MAC_60_14);
	MAC_60_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_15, data_out=>output_MAC_60_15);
	MAC_60_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_16, data_out=>output_MAC_60_16);
	MAC_60_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_17, data_out=>output_MAC_60_17);
	MAC_60_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_18, data_out=>output_MAC_60_18);
	MAC_60_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_19, data_out=>output_MAC_60_19);
	MAC_60_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_20, data_out=>output_MAC_60_20);
	MAC_60_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_21, data_out=>output_MAC_60_21);
	MAC_60_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_22, data_out=>output_MAC_60_22);
	MAC_60_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_23, data_out=>output_MAC_60_23);
	MAC_60_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_24, data_out=>output_MAC_60_24);
	MAC_60_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_25, data_out=>output_MAC_60_25);
	MAC_60_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_26, data_out=>output_MAC_60_26);
	MAC_60_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_27, data_out=>output_MAC_60_27);
	MAC_60_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_28, data_out=>output_MAC_60_28);
	MAC_60_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_29, data_out=>output_MAC_60_29);
	MAC_60_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_30, data_out=>output_MAC_60_30);
	MAC_60_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_31, data_out=>output_MAC_60_31);
	MAC_61_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_0, data_out=>output_MAC_61_0);
	MAC_61_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_1, data_out=>output_MAC_61_1);
	MAC_61_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_2, data_out=>output_MAC_61_2);
	MAC_61_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_3, data_out=>output_MAC_61_3);
	MAC_61_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_4, data_out=>output_MAC_61_4);
	MAC_61_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_5, data_out=>output_MAC_61_5);
	MAC_61_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_6, data_out=>output_MAC_61_6);
	MAC_61_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_7, data_out=>output_MAC_61_7);
	MAC_61_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_8, data_out=>output_MAC_61_8);
	MAC_61_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_9, data_out=>output_MAC_61_9);
	MAC_61_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_10, data_out=>output_MAC_61_10);
	MAC_61_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_11, data_out=>output_MAC_61_11);
	MAC_61_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_12, data_out=>output_MAC_61_12);
	MAC_61_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_13, data_out=>output_MAC_61_13);
	MAC_61_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_14, data_out=>output_MAC_61_14);
	MAC_61_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_15, data_out=>output_MAC_61_15);
	MAC_61_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_16, data_out=>output_MAC_61_16);
	MAC_61_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_17, data_out=>output_MAC_61_17);
	MAC_61_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_18, data_out=>output_MAC_61_18);
	MAC_61_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_19, data_out=>output_MAC_61_19);
	MAC_61_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_20, data_out=>output_MAC_61_20);
	MAC_61_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_21, data_out=>output_MAC_61_21);
	MAC_61_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_22, data_out=>output_MAC_61_22);
	MAC_61_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_23, data_out=>output_MAC_61_23);
	MAC_61_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_24, data_out=>output_MAC_61_24);
	MAC_61_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_25, data_out=>output_MAC_61_25);
	MAC_61_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_26, data_out=>output_MAC_61_26);
	MAC_61_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_27, data_out=>output_MAC_61_27);
	MAC_61_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_28, data_out=>output_MAC_61_28);
	MAC_61_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_29, data_out=>output_MAC_61_29);
	MAC_61_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_30, data_out=>output_MAC_61_30);
	MAC_61_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_31, data_out=>output_MAC_61_31);
	MAC_62_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_0, data_out=>output_MAC_62_0);
	MAC_62_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_1, data_out=>output_MAC_62_1);
	MAC_62_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_2, data_out=>output_MAC_62_2);
	MAC_62_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_3, data_out=>output_MAC_62_3);
	MAC_62_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_4, data_out=>output_MAC_62_4);
	MAC_62_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_5, data_out=>output_MAC_62_5);
	MAC_62_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_6, data_out=>output_MAC_62_6);
	MAC_62_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_7, data_out=>output_MAC_62_7);
	MAC_62_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_8, data_out=>output_MAC_62_8);
	MAC_62_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_9, data_out=>output_MAC_62_9);
	MAC_62_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_10, data_out=>output_MAC_62_10);
	MAC_62_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_11, data_out=>output_MAC_62_11);
	MAC_62_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_12, data_out=>output_MAC_62_12);
	MAC_62_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_13, data_out=>output_MAC_62_13);
	MAC_62_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_14, data_out=>output_MAC_62_14);
	MAC_62_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_15, data_out=>output_MAC_62_15);
	MAC_62_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_16, data_out=>output_MAC_62_16);
	MAC_62_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_17, data_out=>output_MAC_62_17);
	MAC_62_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_18, data_out=>output_MAC_62_18);
	MAC_62_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_19, data_out=>output_MAC_62_19);
	MAC_62_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_20, data_out=>output_MAC_62_20);
	MAC_62_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_21, data_out=>output_MAC_62_21);
	MAC_62_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_22, data_out=>output_MAC_62_22);
	MAC_62_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_23, data_out=>output_MAC_62_23);
	MAC_62_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_24, data_out=>output_MAC_62_24);
	MAC_62_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_25, data_out=>output_MAC_62_25);
	MAC_62_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_26, data_out=>output_MAC_62_26);
	MAC_62_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_27, data_out=>output_MAC_62_27);
	MAC_62_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_28, data_out=>output_MAC_62_28);
	MAC_62_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_29, data_out=>output_MAC_62_29);
	MAC_62_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_30, data_out=>output_MAC_62_30);
	MAC_62_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_31, data_out=>output_MAC_62_31);
	MAC_63_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_0, data_out=>output_MAC_63_0);
	MAC_63_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_1, data_out=>output_MAC_63_1);
	MAC_63_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_2, data_out=>output_MAC_63_2);
	MAC_63_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_3, data_out=>output_MAC_63_3);
	MAC_63_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_4, data_out=>output_MAC_63_4);
	MAC_63_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_5, data_out=>output_MAC_63_5);
	MAC_63_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_6, data_out=>output_MAC_63_6);
	MAC_63_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_7, data_out=>output_MAC_63_7);
	MAC_63_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_8, data_out=>output_MAC_63_8);
	MAC_63_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_9, data_out=>output_MAC_63_9);
	MAC_63_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_10, data_out=>output_MAC_63_10);
	MAC_63_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_11, data_out=>output_MAC_63_11);
	MAC_63_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_12, data_out=>output_MAC_63_12);
	MAC_63_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_13, data_out=>output_MAC_63_13);
	MAC_63_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_14, data_out=>output_MAC_63_14);
	MAC_63_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_15, data_out=>output_MAC_63_15);
	MAC_63_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_16, data_out=>output_MAC_63_16);
	MAC_63_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_17, data_out=>output_MAC_63_17);
	MAC_63_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_18, data_out=>output_MAC_63_18);
	MAC_63_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_19, data_out=>output_MAC_63_19);
	MAC_63_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_20, data_out=>output_MAC_63_20);
	MAC_63_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_21, data_out=>output_MAC_63_21);
	MAC_63_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_22, data_out=>output_MAC_63_22);
	MAC_63_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_23, data_out=>output_MAC_63_23);
	MAC_63_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_24, data_out=>output_MAC_63_24);
	MAC_63_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_25, data_out=>output_MAC_63_25);
	MAC_63_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_26, data_out=>output_MAC_63_26);
	MAC_63_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_27, data_out=>output_MAC_63_27);
	MAC_63_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_28, data_out=>output_MAC_63_28);
	MAC_63_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_29, data_out=>output_MAC_63_29);
	MAC_63_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_30, data_out=>output_MAC_63_30);
	MAC_63_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_31, data_out=>output_MAC_63_31);

	mux_row_0: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_0_0, I1=>output_MAC_0_1, I2=>output_MAC_0_2, I3=>output_MAC_0_3, I4=>output_MAC_0_4, I5=>output_MAC_0_5, I6=>output_MAC_0_6, I7=>output_MAC_0_7, I8=>output_MAC_0_8, I9=>output_MAC_0_9, I10=>output_MAC_0_10, I11=>output_MAC_0_11, I12=>output_MAC_0_12, I13=>output_MAC_0_13, I14=>output_MAC_0_14, I15=>output_MAC_0_15, I16=>output_MAC_0_16, I17=>output_MAC_0_17, I18=>output_MAC_0_18, I19=>output_MAC_0_19, I20=>output_MAC_0_20, I21=>output_MAC_0_21, I22=>output_MAC_0_22, I23=>output_MAC_0_23, I24=>output_MAC_0_24, I25=>output_MAC_0_25, I26=>output_MAC_0_26, I27=>output_MAC_0_27, I28=>output_MAC_0_28, I29=>output_MAC_0_29, I30=>output_MAC_0_30, I31=>output_MAC_0_31, 
		SEL_mux=>SEL_mux, O=>output_row_0);

	mux_row_1: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_1_0, I1=>output_MAC_1_1, I2=>output_MAC_1_2, I3=>output_MAC_1_3, I4=>output_MAC_1_4, I5=>output_MAC_1_5, I6=>output_MAC_1_6, I7=>output_MAC_1_7, I8=>output_MAC_1_8, I9=>output_MAC_1_9, I10=>output_MAC_1_10, I11=>output_MAC_1_11, I12=>output_MAC_1_12, I13=>output_MAC_1_13, I14=>output_MAC_1_14, I15=>output_MAC_1_15, I16=>output_MAC_1_16, I17=>output_MAC_1_17, I18=>output_MAC_1_18, I19=>output_MAC_1_19, I20=>output_MAC_1_20, I21=>output_MAC_1_21, I22=>output_MAC_1_22, I23=>output_MAC_1_23, I24=>output_MAC_1_24, I25=>output_MAC_1_25, I26=>output_MAC_1_26, I27=>output_MAC_1_27, I28=>output_MAC_1_28, I29=>output_MAC_1_29, I30=>output_MAC_1_30, I31=>output_MAC_1_31, 
		SEL_mux=>SEL_mux, O=>output_row_1);

	mux_row_2: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_2_0, I1=>output_MAC_2_1, I2=>output_MAC_2_2, I3=>output_MAC_2_3, I4=>output_MAC_2_4, I5=>output_MAC_2_5, I6=>output_MAC_2_6, I7=>output_MAC_2_7, I8=>output_MAC_2_8, I9=>output_MAC_2_9, I10=>output_MAC_2_10, I11=>output_MAC_2_11, I12=>output_MAC_2_12, I13=>output_MAC_2_13, I14=>output_MAC_2_14, I15=>output_MAC_2_15, I16=>output_MAC_2_16, I17=>output_MAC_2_17, I18=>output_MAC_2_18, I19=>output_MAC_2_19, I20=>output_MAC_2_20, I21=>output_MAC_2_21, I22=>output_MAC_2_22, I23=>output_MAC_2_23, I24=>output_MAC_2_24, I25=>output_MAC_2_25, I26=>output_MAC_2_26, I27=>output_MAC_2_27, I28=>output_MAC_2_28, I29=>output_MAC_2_29, I30=>output_MAC_2_30, I31=>output_MAC_2_31, 
		SEL_mux=>SEL_mux, O=>output_row_2);

	mux_row_3: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_3_0, I1=>output_MAC_3_1, I2=>output_MAC_3_2, I3=>output_MAC_3_3, I4=>output_MAC_3_4, I5=>output_MAC_3_5, I6=>output_MAC_3_6, I7=>output_MAC_3_7, I8=>output_MAC_3_8, I9=>output_MAC_3_9, I10=>output_MAC_3_10, I11=>output_MAC_3_11, I12=>output_MAC_3_12, I13=>output_MAC_3_13, I14=>output_MAC_3_14, I15=>output_MAC_3_15, I16=>output_MAC_3_16, I17=>output_MAC_3_17, I18=>output_MAC_3_18, I19=>output_MAC_3_19, I20=>output_MAC_3_20, I21=>output_MAC_3_21, I22=>output_MAC_3_22, I23=>output_MAC_3_23, I24=>output_MAC_3_24, I25=>output_MAC_3_25, I26=>output_MAC_3_26, I27=>output_MAC_3_27, I28=>output_MAC_3_28, I29=>output_MAC_3_29, I30=>output_MAC_3_30, I31=>output_MAC_3_31, 
		SEL_mux=>SEL_mux, O=>output_row_3);

	mux_row_4: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_4_0, I1=>output_MAC_4_1, I2=>output_MAC_4_2, I3=>output_MAC_4_3, I4=>output_MAC_4_4, I5=>output_MAC_4_5, I6=>output_MAC_4_6, I7=>output_MAC_4_7, I8=>output_MAC_4_8, I9=>output_MAC_4_9, I10=>output_MAC_4_10, I11=>output_MAC_4_11, I12=>output_MAC_4_12, I13=>output_MAC_4_13, I14=>output_MAC_4_14, I15=>output_MAC_4_15, I16=>output_MAC_4_16, I17=>output_MAC_4_17, I18=>output_MAC_4_18, I19=>output_MAC_4_19, I20=>output_MAC_4_20, I21=>output_MAC_4_21, I22=>output_MAC_4_22, I23=>output_MAC_4_23, I24=>output_MAC_4_24, I25=>output_MAC_4_25, I26=>output_MAC_4_26, I27=>output_MAC_4_27, I28=>output_MAC_4_28, I29=>output_MAC_4_29, I30=>output_MAC_4_30, I31=>output_MAC_4_31, 
		SEL_mux=>SEL_mux, O=>output_row_4);

	mux_row_5: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_5_0, I1=>output_MAC_5_1, I2=>output_MAC_5_2, I3=>output_MAC_5_3, I4=>output_MAC_5_4, I5=>output_MAC_5_5, I6=>output_MAC_5_6, I7=>output_MAC_5_7, I8=>output_MAC_5_8, I9=>output_MAC_5_9, I10=>output_MAC_5_10, I11=>output_MAC_5_11, I12=>output_MAC_5_12, I13=>output_MAC_5_13, I14=>output_MAC_5_14, I15=>output_MAC_5_15, I16=>output_MAC_5_16, I17=>output_MAC_5_17, I18=>output_MAC_5_18, I19=>output_MAC_5_19, I20=>output_MAC_5_20, I21=>output_MAC_5_21, I22=>output_MAC_5_22, I23=>output_MAC_5_23, I24=>output_MAC_5_24, I25=>output_MAC_5_25, I26=>output_MAC_5_26, I27=>output_MAC_5_27, I28=>output_MAC_5_28, I29=>output_MAC_5_29, I30=>output_MAC_5_30, I31=>output_MAC_5_31, 
		SEL_mux=>SEL_mux, O=>output_row_5);

	mux_row_6: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_6_0, I1=>output_MAC_6_1, I2=>output_MAC_6_2, I3=>output_MAC_6_3, I4=>output_MAC_6_4, I5=>output_MAC_6_5, I6=>output_MAC_6_6, I7=>output_MAC_6_7, I8=>output_MAC_6_8, I9=>output_MAC_6_9, I10=>output_MAC_6_10, I11=>output_MAC_6_11, I12=>output_MAC_6_12, I13=>output_MAC_6_13, I14=>output_MAC_6_14, I15=>output_MAC_6_15, I16=>output_MAC_6_16, I17=>output_MAC_6_17, I18=>output_MAC_6_18, I19=>output_MAC_6_19, I20=>output_MAC_6_20, I21=>output_MAC_6_21, I22=>output_MAC_6_22, I23=>output_MAC_6_23, I24=>output_MAC_6_24, I25=>output_MAC_6_25, I26=>output_MAC_6_26, I27=>output_MAC_6_27, I28=>output_MAC_6_28, I29=>output_MAC_6_29, I30=>output_MAC_6_30, I31=>output_MAC_6_31, 
		SEL_mux=>SEL_mux, O=>output_row_6);

	mux_row_7: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_7_0, I1=>output_MAC_7_1, I2=>output_MAC_7_2, I3=>output_MAC_7_3, I4=>output_MAC_7_4, I5=>output_MAC_7_5, I6=>output_MAC_7_6, I7=>output_MAC_7_7, I8=>output_MAC_7_8, I9=>output_MAC_7_9, I10=>output_MAC_7_10, I11=>output_MAC_7_11, I12=>output_MAC_7_12, I13=>output_MAC_7_13, I14=>output_MAC_7_14, I15=>output_MAC_7_15, I16=>output_MAC_7_16, I17=>output_MAC_7_17, I18=>output_MAC_7_18, I19=>output_MAC_7_19, I20=>output_MAC_7_20, I21=>output_MAC_7_21, I22=>output_MAC_7_22, I23=>output_MAC_7_23, I24=>output_MAC_7_24, I25=>output_MAC_7_25, I26=>output_MAC_7_26, I27=>output_MAC_7_27, I28=>output_MAC_7_28, I29=>output_MAC_7_29, I30=>output_MAC_7_30, I31=>output_MAC_7_31, 
		SEL_mux=>SEL_mux, O=>output_row_7);

	mux_row_8: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_8_0, I1=>output_MAC_8_1, I2=>output_MAC_8_2, I3=>output_MAC_8_3, I4=>output_MAC_8_4, I5=>output_MAC_8_5, I6=>output_MAC_8_6, I7=>output_MAC_8_7, I8=>output_MAC_8_8, I9=>output_MAC_8_9, I10=>output_MAC_8_10, I11=>output_MAC_8_11, I12=>output_MAC_8_12, I13=>output_MAC_8_13, I14=>output_MAC_8_14, I15=>output_MAC_8_15, I16=>output_MAC_8_16, I17=>output_MAC_8_17, I18=>output_MAC_8_18, I19=>output_MAC_8_19, I20=>output_MAC_8_20, I21=>output_MAC_8_21, I22=>output_MAC_8_22, I23=>output_MAC_8_23, I24=>output_MAC_8_24, I25=>output_MAC_8_25, I26=>output_MAC_8_26, I27=>output_MAC_8_27, I28=>output_MAC_8_28, I29=>output_MAC_8_29, I30=>output_MAC_8_30, I31=>output_MAC_8_31, 
		SEL_mux=>SEL_mux, O=>output_row_8);

	mux_row_9: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_9_0, I1=>output_MAC_9_1, I2=>output_MAC_9_2, I3=>output_MAC_9_3, I4=>output_MAC_9_4, I5=>output_MAC_9_5, I6=>output_MAC_9_6, I7=>output_MAC_9_7, I8=>output_MAC_9_8, I9=>output_MAC_9_9, I10=>output_MAC_9_10, I11=>output_MAC_9_11, I12=>output_MAC_9_12, I13=>output_MAC_9_13, I14=>output_MAC_9_14, I15=>output_MAC_9_15, I16=>output_MAC_9_16, I17=>output_MAC_9_17, I18=>output_MAC_9_18, I19=>output_MAC_9_19, I20=>output_MAC_9_20, I21=>output_MAC_9_21, I22=>output_MAC_9_22, I23=>output_MAC_9_23, I24=>output_MAC_9_24, I25=>output_MAC_9_25, I26=>output_MAC_9_26, I27=>output_MAC_9_27, I28=>output_MAC_9_28, I29=>output_MAC_9_29, I30=>output_MAC_9_30, I31=>output_MAC_9_31, 
		SEL_mux=>SEL_mux, O=>output_row_9);

	mux_row_10: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_10_0, I1=>output_MAC_10_1, I2=>output_MAC_10_2, I3=>output_MAC_10_3, I4=>output_MAC_10_4, I5=>output_MAC_10_5, I6=>output_MAC_10_6, I7=>output_MAC_10_7, I8=>output_MAC_10_8, I9=>output_MAC_10_9, I10=>output_MAC_10_10, I11=>output_MAC_10_11, I12=>output_MAC_10_12, I13=>output_MAC_10_13, I14=>output_MAC_10_14, I15=>output_MAC_10_15, I16=>output_MAC_10_16, I17=>output_MAC_10_17, I18=>output_MAC_10_18, I19=>output_MAC_10_19, I20=>output_MAC_10_20, I21=>output_MAC_10_21, I22=>output_MAC_10_22, I23=>output_MAC_10_23, I24=>output_MAC_10_24, I25=>output_MAC_10_25, I26=>output_MAC_10_26, I27=>output_MAC_10_27, I28=>output_MAC_10_28, I29=>output_MAC_10_29, I30=>output_MAC_10_30, I31=>output_MAC_10_31, 
		SEL_mux=>SEL_mux, O=>output_row_10);

	mux_row_11: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_11_0, I1=>output_MAC_11_1, I2=>output_MAC_11_2, I3=>output_MAC_11_3, I4=>output_MAC_11_4, I5=>output_MAC_11_5, I6=>output_MAC_11_6, I7=>output_MAC_11_7, I8=>output_MAC_11_8, I9=>output_MAC_11_9, I10=>output_MAC_11_10, I11=>output_MAC_11_11, I12=>output_MAC_11_12, I13=>output_MAC_11_13, I14=>output_MAC_11_14, I15=>output_MAC_11_15, I16=>output_MAC_11_16, I17=>output_MAC_11_17, I18=>output_MAC_11_18, I19=>output_MAC_11_19, I20=>output_MAC_11_20, I21=>output_MAC_11_21, I22=>output_MAC_11_22, I23=>output_MAC_11_23, I24=>output_MAC_11_24, I25=>output_MAC_11_25, I26=>output_MAC_11_26, I27=>output_MAC_11_27, I28=>output_MAC_11_28, I29=>output_MAC_11_29, I30=>output_MAC_11_30, I31=>output_MAC_11_31, 
		SEL_mux=>SEL_mux, O=>output_row_11);

	mux_row_12: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_12_0, I1=>output_MAC_12_1, I2=>output_MAC_12_2, I3=>output_MAC_12_3, I4=>output_MAC_12_4, I5=>output_MAC_12_5, I6=>output_MAC_12_6, I7=>output_MAC_12_7, I8=>output_MAC_12_8, I9=>output_MAC_12_9, I10=>output_MAC_12_10, I11=>output_MAC_12_11, I12=>output_MAC_12_12, I13=>output_MAC_12_13, I14=>output_MAC_12_14, I15=>output_MAC_12_15, I16=>output_MAC_12_16, I17=>output_MAC_12_17, I18=>output_MAC_12_18, I19=>output_MAC_12_19, I20=>output_MAC_12_20, I21=>output_MAC_12_21, I22=>output_MAC_12_22, I23=>output_MAC_12_23, I24=>output_MAC_12_24, I25=>output_MAC_12_25, I26=>output_MAC_12_26, I27=>output_MAC_12_27, I28=>output_MAC_12_28, I29=>output_MAC_12_29, I30=>output_MAC_12_30, I31=>output_MAC_12_31, 
		SEL_mux=>SEL_mux, O=>output_row_12);

	mux_row_13: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_13_0, I1=>output_MAC_13_1, I2=>output_MAC_13_2, I3=>output_MAC_13_3, I4=>output_MAC_13_4, I5=>output_MAC_13_5, I6=>output_MAC_13_6, I7=>output_MAC_13_7, I8=>output_MAC_13_8, I9=>output_MAC_13_9, I10=>output_MAC_13_10, I11=>output_MAC_13_11, I12=>output_MAC_13_12, I13=>output_MAC_13_13, I14=>output_MAC_13_14, I15=>output_MAC_13_15, I16=>output_MAC_13_16, I17=>output_MAC_13_17, I18=>output_MAC_13_18, I19=>output_MAC_13_19, I20=>output_MAC_13_20, I21=>output_MAC_13_21, I22=>output_MAC_13_22, I23=>output_MAC_13_23, I24=>output_MAC_13_24, I25=>output_MAC_13_25, I26=>output_MAC_13_26, I27=>output_MAC_13_27, I28=>output_MAC_13_28, I29=>output_MAC_13_29, I30=>output_MAC_13_30, I31=>output_MAC_13_31, 
		SEL_mux=>SEL_mux, O=>output_row_13);

	mux_row_14: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_14_0, I1=>output_MAC_14_1, I2=>output_MAC_14_2, I3=>output_MAC_14_3, I4=>output_MAC_14_4, I5=>output_MAC_14_5, I6=>output_MAC_14_6, I7=>output_MAC_14_7, I8=>output_MAC_14_8, I9=>output_MAC_14_9, I10=>output_MAC_14_10, I11=>output_MAC_14_11, I12=>output_MAC_14_12, I13=>output_MAC_14_13, I14=>output_MAC_14_14, I15=>output_MAC_14_15, I16=>output_MAC_14_16, I17=>output_MAC_14_17, I18=>output_MAC_14_18, I19=>output_MAC_14_19, I20=>output_MAC_14_20, I21=>output_MAC_14_21, I22=>output_MAC_14_22, I23=>output_MAC_14_23, I24=>output_MAC_14_24, I25=>output_MAC_14_25, I26=>output_MAC_14_26, I27=>output_MAC_14_27, I28=>output_MAC_14_28, I29=>output_MAC_14_29, I30=>output_MAC_14_30, I31=>output_MAC_14_31, 
		SEL_mux=>SEL_mux, O=>output_row_14);

	mux_row_15: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_15_0, I1=>output_MAC_15_1, I2=>output_MAC_15_2, I3=>output_MAC_15_3, I4=>output_MAC_15_4, I5=>output_MAC_15_5, I6=>output_MAC_15_6, I7=>output_MAC_15_7, I8=>output_MAC_15_8, I9=>output_MAC_15_9, I10=>output_MAC_15_10, I11=>output_MAC_15_11, I12=>output_MAC_15_12, I13=>output_MAC_15_13, I14=>output_MAC_15_14, I15=>output_MAC_15_15, I16=>output_MAC_15_16, I17=>output_MAC_15_17, I18=>output_MAC_15_18, I19=>output_MAC_15_19, I20=>output_MAC_15_20, I21=>output_MAC_15_21, I22=>output_MAC_15_22, I23=>output_MAC_15_23, I24=>output_MAC_15_24, I25=>output_MAC_15_25, I26=>output_MAC_15_26, I27=>output_MAC_15_27, I28=>output_MAC_15_28, I29=>output_MAC_15_29, I30=>output_MAC_15_30, I31=>output_MAC_15_31, 
		SEL_mux=>SEL_mux, O=>output_row_15);

	mux_row_16: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_16_0, I1=>output_MAC_16_1, I2=>output_MAC_16_2, I3=>output_MAC_16_3, I4=>output_MAC_16_4, I5=>output_MAC_16_5, I6=>output_MAC_16_6, I7=>output_MAC_16_7, I8=>output_MAC_16_8, I9=>output_MAC_16_9, I10=>output_MAC_16_10, I11=>output_MAC_16_11, I12=>output_MAC_16_12, I13=>output_MAC_16_13, I14=>output_MAC_16_14, I15=>output_MAC_16_15, I16=>output_MAC_16_16, I17=>output_MAC_16_17, I18=>output_MAC_16_18, I19=>output_MAC_16_19, I20=>output_MAC_16_20, I21=>output_MAC_16_21, I22=>output_MAC_16_22, I23=>output_MAC_16_23, I24=>output_MAC_16_24, I25=>output_MAC_16_25, I26=>output_MAC_16_26, I27=>output_MAC_16_27, I28=>output_MAC_16_28, I29=>output_MAC_16_29, I30=>output_MAC_16_30, I31=>output_MAC_16_31, 
		SEL_mux=>SEL_mux, O=>output_row_16);

	mux_row_17: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_17_0, I1=>output_MAC_17_1, I2=>output_MAC_17_2, I3=>output_MAC_17_3, I4=>output_MAC_17_4, I5=>output_MAC_17_5, I6=>output_MAC_17_6, I7=>output_MAC_17_7, I8=>output_MAC_17_8, I9=>output_MAC_17_9, I10=>output_MAC_17_10, I11=>output_MAC_17_11, I12=>output_MAC_17_12, I13=>output_MAC_17_13, I14=>output_MAC_17_14, I15=>output_MAC_17_15, I16=>output_MAC_17_16, I17=>output_MAC_17_17, I18=>output_MAC_17_18, I19=>output_MAC_17_19, I20=>output_MAC_17_20, I21=>output_MAC_17_21, I22=>output_MAC_17_22, I23=>output_MAC_17_23, I24=>output_MAC_17_24, I25=>output_MAC_17_25, I26=>output_MAC_17_26, I27=>output_MAC_17_27, I28=>output_MAC_17_28, I29=>output_MAC_17_29, I30=>output_MAC_17_30, I31=>output_MAC_17_31, 
		SEL_mux=>SEL_mux, O=>output_row_17);

	mux_row_18: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_18_0, I1=>output_MAC_18_1, I2=>output_MAC_18_2, I3=>output_MAC_18_3, I4=>output_MAC_18_4, I5=>output_MAC_18_5, I6=>output_MAC_18_6, I7=>output_MAC_18_7, I8=>output_MAC_18_8, I9=>output_MAC_18_9, I10=>output_MAC_18_10, I11=>output_MAC_18_11, I12=>output_MAC_18_12, I13=>output_MAC_18_13, I14=>output_MAC_18_14, I15=>output_MAC_18_15, I16=>output_MAC_18_16, I17=>output_MAC_18_17, I18=>output_MAC_18_18, I19=>output_MAC_18_19, I20=>output_MAC_18_20, I21=>output_MAC_18_21, I22=>output_MAC_18_22, I23=>output_MAC_18_23, I24=>output_MAC_18_24, I25=>output_MAC_18_25, I26=>output_MAC_18_26, I27=>output_MAC_18_27, I28=>output_MAC_18_28, I29=>output_MAC_18_29, I30=>output_MAC_18_30, I31=>output_MAC_18_31, 
		SEL_mux=>SEL_mux, O=>output_row_18);

	mux_row_19: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_19_0, I1=>output_MAC_19_1, I2=>output_MAC_19_2, I3=>output_MAC_19_3, I4=>output_MAC_19_4, I5=>output_MAC_19_5, I6=>output_MAC_19_6, I7=>output_MAC_19_7, I8=>output_MAC_19_8, I9=>output_MAC_19_9, I10=>output_MAC_19_10, I11=>output_MAC_19_11, I12=>output_MAC_19_12, I13=>output_MAC_19_13, I14=>output_MAC_19_14, I15=>output_MAC_19_15, I16=>output_MAC_19_16, I17=>output_MAC_19_17, I18=>output_MAC_19_18, I19=>output_MAC_19_19, I20=>output_MAC_19_20, I21=>output_MAC_19_21, I22=>output_MAC_19_22, I23=>output_MAC_19_23, I24=>output_MAC_19_24, I25=>output_MAC_19_25, I26=>output_MAC_19_26, I27=>output_MAC_19_27, I28=>output_MAC_19_28, I29=>output_MAC_19_29, I30=>output_MAC_19_30, I31=>output_MAC_19_31, 
		SEL_mux=>SEL_mux, O=>output_row_19);

	mux_row_20: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_20_0, I1=>output_MAC_20_1, I2=>output_MAC_20_2, I3=>output_MAC_20_3, I4=>output_MAC_20_4, I5=>output_MAC_20_5, I6=>output_MAC_20_6, I7=>output_MAC_20_7, I8=>output_MAC_20_8, I9=>output_MAC_20_9, I10=>output_MAC_20_10, I11=>output_MAC_20_11, I12=>output_MAC_20_12, I13=>output_MAC_20_13, I14=>output_MAC_20_14, I15=>output_MAC_20_15, I16=>output_MAC_20_16, I17=>output_MAC_20_17, I18=>output_MAC_20_18, I19=>output_MAC_20_19, I20=>output_MAC_20_20, I21=>output_MAC_20_21, I22=>output_MAC_20_22, I23=>output_MAC_20_23, I24=>output_MAC_20_24, I25=>output_MAC_20_25, I26=>output_MAC_20_26, I27=>output_MAC_20_27, I28=>output_MAC_20_28, I29=>output_MAC_20_29, I30=>output_MAC_20_30, I31=>output_MAC_20_31, 
		SEL_mux=>SEL_mux, O=>output_row_20);

	mux_row_21: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_21_0, I1=>output_MAC_21_1, I2=>output_MAC_21_2, I3=>output_MAC_21_3, I4=>output_MAC_21_4, I5=>output_MAC_21_5, I6=>output_MAC_21_6, I7=>output_MAC_21_7, I8=>output_MAC_21_8, I9=>output_MAC_21_9, I10=>output_MAC_21_10, I11=>output_MAC_21_11, I12=>output_MAC_21_12, I13=>output_MAC_21_13, I14=>output_MAC_21_14, I15=>output_MAC_21_15, I16=>output_MAC_21_16, I17=>output_MAC_21_17, I18=>output_MAC_21_18, I19=>output_MAC_21_19, I20=>output_MAC_21_20, I21=>output_MAC_21_21, I22=>output_MAC_21_22, I23=>output_MAC_21_23, I24=>output_MAC_21_24, I25=>output_MAC_21_25, I26=>output_MAC_21_26, I27=>output_MAC_21_27, I28=>output_MAC_21_28, I29=>output_MAC_21_29, I30=>output_MAC_21_30, I31=>output_MAC_21_31, 
		SEL_mux=>SEL_mux, O=>output_row_21);

	mux_row_22: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_22_0, I1=>output_MAC_22_1, I2=>output_MAC_22_2, I3=>output_MAC_22_3, I4=>output_MAC_22_4, I5=>output_MAC_22_5, I6=>output_MAC_22_6, I7=>output_MAC_22_7, I8=>output_MAC_22_8, I9=>output_MAC_22_9, I10=>output_MAC_22_10, I11=>output_MAC_22_11, I12=>output_MAC_22_12, I13=>output_MAC_22_13, I14=>output_MAC_22_14, I15=>output_MAC_22_15, I16=>output_MAC_22_16, I17=>output_MAC_22_17, I18=>output_MAC_22_18, I19=>output_MAC_22_19, I20=>output_MAC_22_20, I21=>output_MAC_22_21, I22=>output_MAC_22_22, I23=>output_MAC_22_23, I24=>output_MAC_22_24, I25=>output_MAC_22_25, I26=>output_MAC_22_26, I27=>output_MAC_22_27, I28=>output_MAC_22_28, I29=>output_MAC_22_29, I30=>output_MAC_22_30, I31=>output_MAC_22_31, 
		SEL_mux=>SEL_mux, O=>output_row_22);

	mux_row_23: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_23_0, I1=>output_MAC_23_1, I2=>output_MAC_23_2, I3=>output_MAC_23_3, I4=>output_MAC_23_4, I5=>output_MAC_23_5, I6=>output_MAC_23_6, I7=>output_MAC_23_7, I8=>output_MAC_23_8, I9=>output_MAC_23_9, I10=>output_MAC_23_10, I11=>output_MAC_23_11, I12=>output_MAC_23_12, I13=>output_MAC_23_13, I14=>output_MAC_23_14, I15=>output_MAC_23_15, I16=>output_MAC_23_16, I17=>output_MAC_23_17, I18=>output_MAC_23_18, I19=>output_MAC_23_19, I20=>output_MAC_23_20, I21=>output_MAC_23_21, I22=>output_MAC_23_22, I23=>output_MAC_23_23, I24=>output_MAC_23_24, I25=>output_MAC_23_25, I26=>output_MAC_23_26, I27=>output_MAC_23_27, I28=>output_MAC_23_28, I29=>output_MAC_23_29, I30=>output_MAC_23_30, I31=>output_MAC_23_31, 
		SEL_mux=>SEL_mux, O=>output_row_23);

	mux_row_24: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_24_0, I1=>output_MAC_24_1, I2=>output_MAC_24_2, I3=>output_MAC_24_3, I4=>output_MAC_24_4, I5=>output_MAC_24_5, I6=>output_MAC_24_6, I7=>output_MAC_24_7, I8=>output_MAC_24_8, I9=>output_MAC_24_9, I10=>output_MAC_24_10, I11=>output_MAC_24_11, I12=>output_MAC_24_12, I13=>output_MAC_24_13, I14=>output_MAC_24_14, I15=>output_MAC_24_15, I16=>output_MAC_24_16, I17=>output_MAC_24_17, I18=>output_MAC_24_18, I19=>output_MAC_24_19, I20=>output_MAC_24_20, I21=>output_MAC_24_21, I22=>output_MAC_24_22, I23=>output_MAC_24_23, I24=>output_MAC_24_24, I25=>output_MAC_24_25, I26=>output_MAC_24_26, I27=>output_MAC_24_27, I28=>output_MAC_24_28, I29=>output_MAC_24_29, I30=>output_MAC_24_30, I31=>output_MAC_24_31, 
		SEL_mux=>SEL_mux, O=>output_row_24);

	mux_row_25: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_25_0, I1=>output_MAC_25_1, I2=>output_MAC_25_2, I3=>output_MAC_25_3, I4=>output_MAC_25_4, I5=>output_MAC_25_5, I6=>output_MAC_25_6, I7=>output_MAC_25_7, I8=>output_MAC_25_8, I9=>output_MAC_25_9, I10=>output_MAC_25_10, I11=>output_MAC_25_11, I12=>output_MAC_25_12, I13=>output_MAC_25_13, I14=>output_MAC_25_14, I15=>output_MAC_25_15, I16=>output_MAC_25_16, I17=>output_MAC_25_17, I18=>output_MAC_25_18, I19=>output_MAC_25_19, I20=>output_MAC_25_20, I21=>output_MAC_25_21, I22=>output_MAC_25_22, I23=>output_MAC_25_23, I24=>output_MAC_25_24, I25=>output_MAC_25_25, I26=>output_MAC_25_26, I27=>output_MAC_25_27, I28=>output_MAC_25_28, I29=>output_MAC_25_29, I30=>output_MAC_25_30, I31=>output_MAC_25_31, 
		SEL_mux=>SEL_mux, O=>output_row_25);

	mux_row_26: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_26_0, I1=>output_MAC_26_1, I2=>output_MAC_26_2, I3=>output_MAC_26_3, I4=>output_MAC_26_4, I5=>output_MAC_26_5, I6=>output_MAC_26_6, I7=>output_MAC_26_7, I8=>output_MAC_26_8, I9=>output_MAC_26_9, I10=>output_MAC_26_10, I11=>output_MAC_26_11, I12=>output_MAC_26_12, I13=>output_MAC_26_13, I14=>output_MAC_26_14, I15=>output_MAC_26_15, I16=>output_MAC_26_16, I17=>output_MAC_26_17, I18=>output_MAC_26_18, I19=>output_MAC_26_19, I20=>output_MAC_26_20, I21=>output_MAC_26_21, I22=>output_MAC_26_22, I23=>output_MAC_26_23, I24=>output_MAC_26_24, I25=>output_MAC_26_25, I26=>output_MAC_26_26, I27=>output_MAC_26_27, I28=>output_MAC_26_28, I29=>output_MAC_26_29, I30=>output_MAC_26_30, I31=>output_MAC_26_31, 
		SEL_mux=>SEL_mux, O=>output_row_26);

	mux_row_27: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_27_0, I1=>output_MAC_27_1, I2=>output_MAC_27_2, I3=>output_MAC_27_3, I4=>output_MAC_27_4, I5=>output_MAC_27_5, I6=>output_MAC_27_6, I7=>output_MAC_27_7, I8=>output_MAC_27_8, I9=>output_MAC_27_9, I10=>output_MAC_27_10, I11=>output_MAC_27_11, I12=>output_MAC_27_12, I13=>output_MAC_27_13, I14=>output_MAC_27_14, I15=>output_MAC_27_15, I16=>output_MAC_27_16, I17=>output_MAC_27_17, I18=>output_MAC_27_18, I19=>output_MAC_27_19, I20=>output_MAC_27_20, I21=>output_MAC_27_21, I22=>output_MAC_27_22, I23=>output_MAC_27_23, I24=>output_MAC_27_24, I25=>output_MAC_27_25, I26=>output_MAC_27_26, I27=>output_MAC_27_27, I28=>output_MAC_27_28, I29=>output_MAC_27_29, I30=>output_MAC_27_30, I31=>output_MAC_27_31, 
		SEL_mux=>SEL_mux, O=>output_row_27);

	mux_row_28: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_28_0, I1=>output_MAC_28_1, I2=>output_MAC_28_2, I3=>output_MAC_28_3, I4=>output_MAC_28_4, I5=>output_MAC_28_5, I6=>output_MAC_28_6, I7=>output_MAC_28_7, I8=>output_MAC_28_8, I9=>output_MAC_28_9, I10=>output_MAC_28_10, I11=>output_MAC_28_11, I12=>output_MAC_28_12, I13=>output_MAC_28_13, I14=>output_MAC_28_14, I15=>output_MAC_28_15, I16=>output_MAC_28_16, I17=>output_MAC_28_17, I18=>output_MAC_28_18, I19=>output_MAC_28_19, I20=>output_MAC_28_20, I21=>output_MAC_28_21, I22=>output_MAC_28_22, I23=>output_MAC_28_23, I24=>output_MAC_28_24, I25=>output_MAC_28_25, I26=>output_MAC_28_26, I27=>output_MAC_28_27, I28=>output_MAC_28_28, I29=>output_MAC_28_29, I30=>output_MAC_28_30, I31=>output_MAC_28_31, 
		SEL_mux=>SEL_mux, O=>output_row_28);

	mux_row_29: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_29_0, I1=>output_MAC_29_1, I2=>output_MAC_29_2, I3=>output_MAC_29_3, I4=>output_MAC_29_4, I5=>output_MAC_29_5, I6=>output_MAC_29_6, I7=>output_MAC_29_7, I8=>output_MAC_29_8, I9=>output_MAC_29_9, I10=>output_MAC_29_10, I11=>output_MAC_29_11, I12=>output_MAC_29_12, I13=>output_MAC_29_13, I14=>output_MAC_29_14, I15=>output_MAC_29_15, I16=>output_MAC_29_16, I17=>output_MAC_29_17, I18=>output_MAC_29_18, I19=>output_MAC_29_19, I20=>output_MAC_29_20, I21=>output_MAC_29_21, I22=>output_MAC_29_22, I23=>output_MAC_29_23, I24=>output_MAC_29_24, I25=>output_MAC_29_25, I26=>output_MAC_29_26, I27=>output_MAC_29_27, I28=>output_MAC_29_28, I29=>output_MAC_29_29, I30=>output_MAC_29_30, I31=>output_MAC_29_31, 
		SEL_mux=>SEL_mux, O=>output_row_29);

	mux_row_30: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_30_0, I1=>output_MAC_30_1, I2=>output_MAC_30_2, I3=>output_MAC_30_3, I4=>output_MAC_30_4, I5=>output_MAC_30_5, I6=>output_MAC_30_6, I7=>output_MAC_30_7, I8=>output_MAC_30_8, I9=>output_MAC_30_9, I10=>output_MAC_30_10, I11=>output_MAC_30_11, I12=>output_MAC_30_12, I13=>output_MAC_30_13, I14=>output_MAC_30_14, I15=>output_MAC_30_15, I16=>output_MAC_30_16, I17=>output_MAC_30_17, I18=>output_MAC_30_18, I19=>output_MAC_30_19, I20=>output_MAC_30_20, I21=>output_MAC_30_21, I22=>output_MAC_30_22, I23=>output_MAC_30_23, I24=>output_MAC_30_24, I25=>output_MAC_30_25, I26=>output_MAC_30_26, I27=>output_MAC_30_27, I28=>output_MAC_30_28, I29=>output_MAC_30_29, I30=>output_MAC_30_30, I31=>output_MAC_30_31, 
		SEL_mux=>SEL_mux, O=>output_row_30);

	mux_row_31: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_31_0, I1=>output_MAC_31_1, I2=>output_MAC_31_2, I3=>output_MAC_31_3, I4=>output_MAC_31_4, I5=>output_MAC_31_5, I6=>output_MAC_31_6, I7=>output_MAC_31_7, I8=>output_MAC_31_8, I9=>output_MAC_31_9, I10=>output_MAC_31_10, I11=>output_MAC_31_11, I12=>output_MAC_31_12, I13=>output_MAC_31_13, I14=>output_MAC_31_14, I15=>output_MAC_31_15, I16=>output_MAC_31_16, I17=>output_MAC_31_17, I18=>output_MAC_31_18, I19=>output_MAC_31_19, I20=>output_MAC_31_20, I21=>output_MAC_31_21, I22=>output_MAC_31_22, I23=>output_MAC_31_23, I24=>output_MAC_31_24, I25=>output_MAC_31_25, I26=>output_MAC_31_26, I27=>output_MAC_31_27, I28=>output_MAC_31_28, I29=>output_MAC_31_29, I30=>output_MAC_31_30, I31=>output_MAC_31_31, 
		SEL_mux=>SEL_mux, O=>output_row_31);

	mux_row_32: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_32_0, I1=>output_MAC_32_1, I2=>output_MAC_32_2, I3=>output_MAC_32_3, I4=>output_MAC_32_4, I5=>output_MAC_32_5, I6=>output_MAC_32_6, I7=>output_MAC_32_7, I8=>output_MAC_32_8, I9=>output_MAC_32_9, I10=>output_MAC_32_10, I11=>output_MAC_32_11, I12=>output_MAC_32_12, I13=>output_MAC_32_13, I14=>output_MAC_32_14, I15=>output_MAC_32_15, I16=>output_MAC_32_16, I17=>output_MAC_32_17, I18=>output_MAC_32_18, I19=>output_MAC_32_19, I20=>output_MAC_32_20, I21=>output_MAC_32_21, I22=>output_MAC_32_22, I23=>output_MAC_32_23, I24=>output_MAC_32_24, I25=>output_MAC_32_25, I26=>output_MAC_32_26, I27=>output_MAC_32_27, I28=>output_MAC_32_28, I29=>output_MAC_32_29, I30=>output_MAC_32_30, I31=>output_MAC_32_31, 
		SEL_mux=>SEL_mux, O=>output_row_32);

	mux_row_33: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_33_0, I1=>output_MAC_33_1, I2=>output_MAC_33_2, I3=>output_MAC_33_3, I4=>output_MAC_33_4, I5=>output_MAC_33_5, I6=>output_MAC_33_6, I7=>output_MAC_33_7, I8=>output_MAC_33_8, I9=>output_MAC_33_9, I10=>output_MAC_33_10, I11=>output_MAC_33_11, I12=>output_MAC_33_12, I13=>output_MAC_33_13, I14=>output_MAC_33_14, I15=>output_MAC_33_15, I16=>output_MAC_33_16, I17=>output_MAC_33_17, I18=>output_MAC_33_18, I19=>output_MAC_33_19, I20=>output_MAC_33_20, I21=>output_MAC_33_21, I22=>output_MAC_33_22, I23=>output_MAC_33_23, I24=>output_MAC_33_24, I25=>output_MAC_33_25, I26=>output_MAC_33_26, I27=>output_MAC_33_27, I28=>output_MAC_33_28, I29=>output_MAC_33_29, I30=>output_MAC_33_30, I31=>output_MAC_33_31, 
		SEL_mux=>SEL_mux, O=>output_row_33);

	mux_row_34: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_34_0, I1=>output_MAC_34_1, I2=>output_MAC_34_2, I3=>output_MAC_34_3, I4=>output_MAC_34_4, I5=>output_MAC_34_5, I6=>output_MAC_34_6, I7=>output_MAC_34_7, I8=>output_MAC_34_8, I9=>output_MAC_34_9, I10=>output_MAC_34_10, I11=>output_MAC_34_11, I12=>output_MAC_34_12, I13=>output_MAC_34_13, I14=>output_MAC_34_14, I15=>output_MAC_34_15, I16=>output_MAC_34_16, I17=>output_MAC_34_17, I18=>output_MAC_34_18, I19=>output_MAC_34_19, I20=>output_MAC_34_20, I21=>output_MAC_34_21, I22=>output_MAC_34_22, I23=>output_MAC_34_23, I24=>output_MAC_34_24, I25=>output_MAC_34_25, I26=>output_MAC_34_26, I27=>output_MAC_34_27, I28=>output_MAC_34_28, I29=>output_MAC_34_29, I30=>output_MAC_34_30, I31=>output_MAC_34_31, 
		SEL_mux=>SEL_mux, O=>output_row_34);

	mux_row_35: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_35_0, I1=>output_MAC_35_1, I2=>output_MAC_35_2, I3=>output_MAC_35_3, I4=>output_MAC_35_4, I5=>output_MAC_35_5, I6=>output_MAC_35_6, I7=>output_MAC_35_7, I8=>output_MAC_35_8, I9=>output_MAC_35_9, I10=>output_MAC_35_10, I11=>output_MAC_35_11, I12=>output_MAC_35_12, I13=>output_MAC_35_13, I14=>output_MAC_35_14, I15=>output_MAC_35_15, I16=>output_MAC_35_16, I17=>output_MAC_35_17, I18=>output_MAC_35_18, I19=>output_MAC_35_19, I20=>output_MAC_35_20, I21=>output_MAC_35_21, I22=>output_MAC_35_22, I23=>output_MAC_35_23, I24=>output_MAC_35_24, I25=>output_MAC_35_25, I26=>output_MAC_35_26, I27=>output_MAC_35_27, I28=>output_MAC_35_28, I29=>output_MAC_35_29, I30=>output_MAC_35_30, I31=>output_MAC_35_31, 
		SEL_mux=>SEL_mux, O=>output_row_35);

	mux_row_36: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_36_0, I1=>output_MAC_36_1, I2=>output_MAC_36_2, I3=>output_MAC_36_3, I4=>output_MAC_36_4, I5=>output_MAC_36_5, I6=>output_MAC_36_6, I7=>output_MAC_36_7, I8=>output_MAC_36_8, I9=>output_MAC_36_9, I10=>output_MAC_36_10, I11=>output_MAC_36_11, I12=>output_MAC_36_12, I13=>output_MAC_36_13, I14=>output_MAC_36_14, I15=>output_MAC_36_15, I16=>output_MAC_36_16, I17=>output_MAC_36_17, I18=>output_MAC_36_18, I19=>output_MAC_36_19, I20=>output_MAC_36_20, I21=>output_MAC_36_21, I22=>output_MAC_36_22, I23=>output_MAC_36_23, I24=>output_MAC_36_24, I25=>output_MAC_36_25, I26=>output_MAC_36_26, I27=>output_MAC_36_27, I28=>output_MAC_36_28, I29=>output_MAC_36_29, I30=>output_MAC_36_30, I31=>output_MAC_36_31, 
		SEL_mux=>SEL_mux, O=>output_row_36);

	mux_row_37: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_37_0, I1=>output_MAC_37_1, I2=>output_MAC_37_2, I3=>output_MAC_37_3, I4=>output_MAC_37_4, I5=>output_MAC_37_5, I6=>output_MAC_37_6, I7=>output_MAC_37_7, I8=>output_MAC_37_8, I9=>output_MAC_37_9, I10=>output_MAC_37_10, I11=>output_MAC_37_11, I12=>output_MAC_37_12, I13=>output_MAC_37_13, I14=>output_MAC_37_14, I15=>output_MAC_37_15, I16=>output_MAC_37_16, I17=>output_MAC_37_17, I18=>output_MAC_37_18, I19=>output_MAC_37_19, I20=>output_MAC_37_20, I21=>output_MAC_37_21, I22=>output_MAC_37_22, I23=>output_MAC_37_23, I24=>output_MAC_37_24, I25=>output_MAC_37_25, I26=>output_MAC_37_26, I27=>output_MAC_37_27, I28=>output_MAC_37_28, I29=>output_MAC_37_29, I30=>output_MAC_37_30, I31=>output_MAC_37_31, 
		SEL_mux=>SEL_mux, O=>output_row_37);

	mux_row_38: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_38_0, I1=>output_MAC_38_1, I2=>output_MAC_38_2, I3=>output_MAC_38_3, I4=>output_MAC_38_4, I5=>output_MAC_38_5, I6=>output_MAC_38_6, I7=>output_MAC_38_7, I8=>output_MAC_38_8, I9=>output_MAC_38_9, I10=>output_MAC_38_10, I11=>output_MAC_38_11, I12=>output_MAC_38_12, I13=>output_MAC_38_13, I14=>output_MAC_38_14, I15=>output_MAC_38_15, I16=>output_MAC_38_16, I17=>output_MAC_38_17, I18=>output_MAC_38_18, I19=>output_MAC_38_19, I20=>output_MAC_38_20, I21=>output_MAC_38_21, I22=>output_MAC_38_22, I23=>output_MAC_38_23, I24=>output_MAC_38_24, I25=>output_MAC_38_25, I26=>output_MAC_38_26, I27=>output_MAC_38_27, I28=>output_MAC_38_28, I29=>output_MAC_38_29, I30=>output_MAC_38_30, I31=>output_MAC_38_31, 
		SEL_mux=>SEL_mux, O=>output_row_38);

	mux_row_39: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_39_0, I1=>output_MAC_39_1, I2=>output_MAC_39_2, I3=>output_MAC_39_3, I4=>output_MAC_39_4, I5=>output_MAC_39_5, I6=>output_MAC_39_6, I7=>output_MAC_39_7, I8=>output_MAC_39_8, I9=>output_MAC_39_9, I10=>output_MAC_39_10, I11=>output_MAC_39_11, I12=>output_MAC_39_12, I13=>output_MAC_39_13, I14=>output_MAC_39_14, I15=>output_MAC_39_15, I16=>output_MAC_39_16, I17=>output_MAC_39_17, I18=>output_MAC_39_18, I19=>output_MAC_39_19, I20=>output_MAC_39_20, I21=>output_MAC_39_21, I22=>output_MAC_39_22, I23=>output_MAC_39_23, I24=>output_MAC_39_24, I25=>output_MAC_39_25, I26=>output_MAC_39_26, I27=>output_MAC_39_27, I28=>output_MAC_39_28, I29=>output_MAC_39_29, I30=>output_MAC_39_30, I31=>output_MAC_39_31, 
		SEL_mux=>SEL_mux, O=>output_row_39);

	mux_row_40: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_40_0, I1=>output_MAC_40_1, I2=>output_MAC_40_2, I3=>output_MAC_40_3, I4=>output_MAC_40_4, I5=>output_MAC_40_5, I6=>output_MAC_40_6, I7=>output_MAC_40_7, I8=>output_MAC_40_8, I9=>output_MAC_40_9, I10=>output_MAC_40_10, I11=>output_MAC_40_11, I12=>output_MAC_40_12, I13=>output_MAC_40_13, I14=>output_MAC_40_14, I15=>output_MAC_40_15, I16=>output_MAC_40_16, I17=>output_MAC_40_17, I18=>output_MAC_40_18, I19=>output_MAC_40_19, I20=>output_MAC_40_20, I21=>output_MAC_40_21, I22=>output_MAC_40_22, I23=>output_MAC_40_23, I24=>output_MAC_40_24, I25=>output_MAC_40_25, I26=>output_MAC_40_26, I27=>output_MAC_40_27, I28=>output_MAC_40_28, I29=>output_MAC_40_29, I30=>output_MAC_40_30, I31=>output_MAC_40_31, 
		SEL_mux=>SEL_mux, O=>output_row_40);

	mux_row_41: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_41_0, I1=>output_MAC_41_1, I2=>output_MAC_41_2, I3=>output_MAC_41_3, I4=>output_MAC_41_4, I5=>output_MAC_41_5, I6=>output_MAC_41_6, I7=>output_MAC_41_7, I8=>output_MAC_41_8, I9=>output_MAC_41_9, I10=>output_MAC_41_10, I11=>output_MAC_41_11, I12=>output_MAC_41_12, I13=>output_MAC_41_13, I14=>output_MAC_41_14, I15=>output_MAC_41_15, I16=>output_MAC_41_16, I17=>output_MAC_41_17, I18=>output_MAC_41_18, I19=>output_MAC_41_19, I20=>output_MAC_41_20, I21=>output_MAC_41_21, I22=>output_MAC_41_22, I23=>output_MAC_41_23, I24=>output_MAC_41_24, I25=>output_MAC_41_25, I26=>output_MAC_41_26, I27=>output_MAC_41_27, I28=>output_MAC_41_28, I29=>output_MAC_41_29, I30=>output_MAC_41_30, I31=>output_MAC_41_31, 
		SEL_mux=>SEL_mux, O=>output_row_41);

	mux_row_42: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_42_0, I1=>output_MAC_42_1, I2=>output_MAC_42_2, I3=>output_MAC_42_3, I4=>output_MAC_42_4, I5=>output_MAC_42_5, I6=>output_MAC_42_6, I7=>output_MAC_42_7, I8=>output_MAC_42_8, I9=>output_MAC_42_9, I10=>output_MAC_42_10, I11=>output_MAC_42_11, I12=>output_MAC_42_12, I13=>output_MAC_42_13, I14=>output_MAC_42_14, I15=>output_MAC_42_15, I16=>output_MAC_42_16, I17=>output_MAC_42_17, I18=>output_MAC_42_18, I19=>output_MAC_42_19, I20=>output_MAC_42_20, I21=>output_MAC_42_21, I22=>output_MAC_42_22, I23=>output_MAC_42_23, I24=>output_MAC_42_24, I25=>output_MAC_42_25, I26=>output_MAC_42_26, I27=>output_MAC_42_27, I28=>output_MAC_42_28, I29=>output_MAC_42_29, I30=>output_MAC_42_30, I31=>output_MAC_42_31, 
		SEL_mux=>SEL_mux, O=>output_row_42);

	mux_row_43: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_43_0, I1=>output_MAC_43_1, I2=>output_MAC_43_2, I3=>output_MAC_43_3, I4=>output_MAC_43_4, I5=>output_MAC_43_5, I6=>output_MAC_43_6, I7=>output_MAC_43_7, I8=>output_MAC_43_8, I9=>output_MAC_43_9, I10=>output_MAC_43_10, I11=>output_MAC_43_11, I12=>output_MAC_43_12, I13=>output_MAC_43_13, I14=>output_MAC_43_14, I15=>output_MAC_43_15, I16=>output_MAC_43_16, I17=>output_MAC_43_17, I18=>output_MAC_43_18, I19=>output_MAC_43_19, I20=>output_MAC_43_20, I21=>output_MAC_43_21, I22=>output_MAC_43_22, I23=>output_MAC_43_23, I24=>output_MAC_43_24, I25=>output_MAC_43_25, I26=>output_MAC_43_26, I27=>output_MAC_43_27, I28=>output_MAC_43_28, I29=>output_MAC_43_29, I30=>output_MAC_43_30, I31=>output_MAC_43_31, 
		SEL_mux=>SEL_mux, O=>output_row_43);

	mux_row_44: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_44_0, I1=>output_MAC_44_1, I2=>output_MAC_44_2, I3=>output_MAC_44_3, I4=>output_MAC_44_4, I5=>output_MAC_44_5, I6=>output_MAC_44_6, I7=>output_MAC_44_7, I8=>output_MAC_44_8, I9=>output_MAC_44_9, I10=>output_MAC_44_10, I11=>output_MAC_44_11, I12=>output_MAC_44_12, I13=>output_MAC_44_13, I14=>output_MAC_44_14, I15=>output_MAC_44_15, I16=>output_MAC_44_16, I17=>output_MAC_44_17, I18=>output_MAC_44_18, I19=>output_MAC_44_19, I20=>output_MAC_44_20, I21=>output_MAC_44_21, I22=>output_MAC_44_22, I23=>output_MAC_44_23, I24=>output_MAC_44_24, I25=>output_MAC_44_25, I26=>output_MAC_44_26, I27=>output_MAC_44_27, I28=>output_MAC_44_28, I29=>output_MAC_44_29, I30=>output_MAC_44_30, I31=>output_MAC_44_31, 
		SEL_mux=>SEL_mux, O=>output_row_44);

	mux_row_45: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_45_0, I1=>output_MAC_45_1, I2=>output_MAC_45_2, I3=>output_MAC_45_3, I4=>output_MAC_45_4, I5=>output_MAC_45_5, I6=>output_MAC_45_6, I7=>output_MAC_45_7, I8=>output_MAC_45_8, I9=>output_MAC_45_9, I10=>output_MAC_45_10, I11=>output_MAC_45_11, I12=>output_MAC_45_12, I13=>output_MAC_45_13, I14=>output_MAC_45_14, I15=>output_MAC_45_15, I16=>output_MAC_45_16, I17=>output_MAC_45_17, I18=>output_MAC_45_18, I19=>output_MAC_45_19, I20=>output_MAC_45_20, I21=>output_MAC_45_21, I22=>output_MAC_45_22, I23=>output_MAC_45_23, I24=>output_MAC_45_24, I25=>output_MAC_45_25, I26=>output_MAC_45_26, I27=>output_MAC_45_27, I28=>output_MAC_45_28, I29=>output_MAC_45_29, I30=>output_MAC_45_30, I31=>output_MAC_45_31, 
		SEL_mux=>SEL_mux, O=>output_row_45);

	mux_row_46: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_46_0, I1=>output_MAC_46_1, I2=>output_MAC_46_2, I3=>output_MAC_46_3, I4=>output_MAC_46_4, I5=>output_MAC_46_5, I6=>output_MAC_46_6, I7=>output_MAC_46_7, I8=>output_MAC_46_8, I9=>output_MAC_46_9, I10=>output_MAC_46_10, I11=>output_MAC_46_11, I12=>output_MAC_46_12, I13=>output_MAC_46_13, I14=>output_MAC_46_14, I15=>output_MAC_46_15, I16=>output_MAC_46_16, I17=>output_MAC_46_17, I18=>output_MAC_46_18, I19=>output_MAC_46_19, I20=>output_MAC_46_20, I21=>output_MAC_46_21, I22=>output_MAC_46_22, I23=>output_MAC_46_23, I24=>output_MAC_46_24, I25=>output_MAC_46_25, I26=>output_MAC_46_26, I27=>output_MAC_46_27, I28=>output_MAC_46_28, I29=>output_MAC_46_29, I30=>output_MAC_46_30, I31=>output_MAC_46_31, 
		SEL_mux=>SEL_mux, O=>output_row_46);

	mux_row_47: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_47_0, I1=>output_MAC_47_1, I2=>output_MAC_47_2, I3=>output_MAC_47_3, I4=>output_MAC_47_4, I5=>output_MAC_47_5, I6=>output_MAC_47_6, I7=>output_MAC_47_7, I8=>output_MAC_47_8, I9=>output_MAC_47_9, I10=>output_MAC_47_10, I11=>output_MAC_47_11, I12=>output_MAC_47_12, I13=>output_MAC_47_13, I14=>output_MAC_47_14, I15=>output_MAC_47_15, I16=>output_MAC_47_16, I17=>output_MAC_47_17, I18=>output_MAC_47_18, I19=>output_MAC_47_19, I20=>output_MAC_47_20, I21=>output_MAC_47_21, I22=>output_MAC_47_22, I23=>output_MAC_47_23, I24=>output_MAC_47_24, I25=>output_MAC_47_25, I26=>output_MAC_47_26, I27=>output_MAC_47_27, I28=>output_MAC_47_28, I29=>output_MAC_47_29, I30=>output_MAC_47_30, I31=>output_MAC_47_31, 
		SEL_mux=>SEL_mux, O=>output_row_47);

	mux_row_48: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_48_0, I1=>output_MAC_48_1, I2=>output_MAC_48_2, I3=>output_MAC_48_3, I4=>output_MAC_48_4, I5=>output_MAC_48_5, I6=>output_MAC_48_6, I7=>output_MAC_48_7, I8=>output_MAC_48_8, I9=>output_MAC_48_9, I10=>output_MAC_48_10, I11=>output_MAC_48_11, I12=>output_MAC_48_12, I13=>output_MAC_48_13, I14=>output_MAC_48_14, I15=>output_MAC_48_15, I16=>output_MAC_48_16, I17=>output_MAC_48_17, I18=>output_MAC_48_18, I19=>output_MAC_48_19, I20=>output_MAC_48_20, I21=>output_MAC_48_21, I22=>output_MAC_48_22, I23=>output_MAC_48_23, I24=>output_MAC_48_24, I25=>output_MAC_48_25, I26=>output_MAC_48_26, I27=>output_MAC_48_27, I28=>output_MAC_48_28, I29=>output_MAC_48_29, I30=>output_MAC_48_30, I31=>output_MAC_48_31, 
		SEL_mux=>SEL_mux, O=>output_row_48);

	mux_row_49: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_49_0, I1=>output_MAC_49_1, I2=>output_MAC_49_2, I3=>output_MAC_49_3, I4=>output_MAC_49_4, I5=>output_MAC_49_5, I6=>output_MAC_49_6, I7=>output_MAC_49_7, I8=>output_MAC_49_8, I9=>output_MAC_49_9, I10=>output_MAC_49_10, I11=>output_MAC_49_11, I12=>output_MAC_49_12, I13=>output_MAC_49_13, I14=>output_MAC_49_14, I15=>output_MAC_49_15, I16=>output_MAC_49_16, I17=>output_MAC_49_17, I18=>output_MAC_49_18, I19=>output_MAC_49_19, I20=>output_MAC_49_20, I21=>output_MAC_49_21, I22=>output_MAC_49_22, I23=>output_MAC_49_23, I24=>output_MAC_49_24, I25=>output_MAC_49_25, I26=>output_MAC_49_26, I27=>output_MAC_49_27, I28=>output_MAC_49_28, I29=>output_MAC_49_29, I30=>output_MAC_49_30, I31=>output_MAC_49_31, 
		SEL_mux=>SEL_mux, O=>output_row_49);

	mux_row_50: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_50_0, I1=>output_MAC_50_1, I2=>output_MAC_50_2, I3=>output_MAC_50_3, I4=>output_MAC_50_4, I5=>output_MAC_50_5, I6=>output_MAC_50_6, I7=>output_MAC_50_7, I8=>output_MAC_50_8, I9=>output_MAC_50_9, I10=>output_MAC_50_10, I11=>output_MAC_50_11, I12=>output_MAC_50_12, I13=>output_MAC_50_13, I14=>output_MAC_50_14, I15=>output_MAC_50_15, I16=>output_MAC_50_16, I17=>output_MAC_50_17, I18=>output_MAC_50_18, I19=>output_MAC_50_19, I20=>output_MAC_50_20, I21=>output_MAC_50_21, I22=>output_MAC_50_22, I23=>output_MAC_50_23, I24=>output_MAC_50_24, I25=>output_MAC_50_25, I26=>output_MAC_50_26, I27=>output_MAC_50_27, I28=>output_MAC_50_28, I29=>output_MAC_50_29, I30=>output_MAC_50_30, I31=>output_MAC_50_31, 
		SEL_mux=>SEL_mux, O=>output_row_50);

	mux_row_51: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_51_0, I1=>output_MAC_51_1, I2=>output_MAC_51_2, I3=>output_MAC_51_3, I4=>output_MAC_51_4, I5=>output_MAC_51_5, I6=>output_MAC_51_6, I7=>output_MAC_51_7, I8=>output_MAC_51_8, I9=>output_MAC_51_9, I10=>output_MAC_51_10, I11=>output_MAC_51_11, I12=>output_MAC_51_12, I13=>output_MAC_51_13, I14=>output_MAC_51_14, I15=>output_MAC_51_15, I16=>output_MAC_51_16, I17=>output_MAC_51_17, I18=>output_MAC_51_18, I19=>output_MAC_51_19, I20=>output_MAC_51_20, I21=>output_MAC_51_21, I22=>output_MAC_51_22, I23=>output_MAC_51_23, I24=>output_MAC_51_24, I25=>output_MAC_51_25, I26=>output_MAC_51_26, I27=>output_MAC_51_27, I28=>output_MAC_51_28, I29=>output_MAC_51_29, I30=>output_MAC_51_30, I31=>output_MAC_51_31, 
		SEL_mux=>SEL_mux, O=>output_row_51);

	mux_row_52: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_52_0, I1=>output_MAC_52_1, I2=>output_MAC_52_2, I3=>output_MAC_52_3, I4=>output_MAC_52_4, I5=>output_MAC_52_5, I6=>output_MAC_52_6, I7=>output_MAC_52_7, I8=>output_MAC_52_8, I9=>output_MAC_52_9, I10=>output_MAC_52_10, I11=>output_MAC_52_11, I12=>output_MAC_52_12, I13=>output_MAC_52_13, I14=>output_MAC_52_14, I15=>output_MAC_52_15, I16=>output_MAC_52_16, I17=>output_MAC_52_17, I18=>output_MAC_52_18, I19=>output_MAC_52_19, I20=>output_MAC_52_20, I21=>output_MAC_52_21, I22=>output_MAC_52_22, I23=>output_MAC_52_23, I24=>output_MAC_52_24, I25=>output_MAC_52_25, I26=>output_MAC_52_26, I27=>output_MAC_52_27, I28=>output_MAC_52_28, I29=>output_MAC_52_29, I30=>output_MAC_52_30, I31=>output_MAC_52_31, 
		SEL_mux=>SEL_mux, O=>output_row_52);

	mux_row_53: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_53_0, I1=>output_MAC_53_1, I2=>output_MAC_53_2, I3=>output_MAC_53_3, I4=>output_MAC_53_4, I5=>output_MAC_53_5, I6=>output_MAC_53_6, I7=>output_MAC_53_7, I8=>output_MAC_53_8, I9=>output_MAC_53_9, I10=>output_MAC_53_10, I11=>output_MAC_53_11, I12=>output_MAC_53_12, I13=>output_MAC_53_13, I14=>output_MAC_53_14, I15=>output_MAC_53_15, I16=>output_MAC_53_16, I17=>output_MAC_53_17, I18=>output_MAC_53_18, I19=>output_MAC_53_19, I20=>output_MAC_53_20, I21=>output_MAC_53_21, I22=>output_MAC_53_22, I23=>output_MAC_53_23, I24=>output_MAC_53_24, I25=>output_MAC_53_25, I26=>output_MAC_53_26, I27=>output_MAC_53_27, I28=>output_MAC_53_28, I29=>output_MAC_53_29, I30=>output_MAC_53_30, I31=>output_MAC_53_31, 
		SEL_mux=>SEL_mux, O=>output_row_53);

	mux_row_54: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_54_0, I1=>output_MAC_54_1, I2=>output_MAC_54_2, I3=>output_MAC_54_3, I4=>output_MAC_54_4, I5=>output_MAC_54_5, I6=>output_MAC_54_6, I7=>output_MAC_54_7, I8=>output_MAC_54_8, I9=>output_MAC_54_9, I10=>output_MAC_54_10, I11=>output_MAC_54_11, I12=>output_MAC_54_12, I13=>output_MAC_54_13, I14=>output_MAC_54_14, I15=>output_MAC_54_15, I16=>output_MAC_54_16, I17=>output_MAC_54_17, I18=>output_MAC_54_18, I19=>output_MAC_54_19, I20=>output_MAC_54_20, I21=>output_MAC_54_21, I22=>output_MAC_54_22, I23=>output_MAC_54_23, I24=>output_MAC_54_24, I25=>output_MAC_54_25, I26=>output_MAC_54_26, I27=>output_MAC_54_27, I28=>output_MAC_54_28, I29=>output_MAC_54_29, I30=>output_MAC_54_30, I31=>output_MAC_54_31, 
		SEL_mux=>SEL_mux, O=>output_row_54);

	mux_row_55: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_55_0, I1=>output_MAC_55_1, I2=>output_MAC_55_2, I3=>output_MAC_55_3, I4=>output_MAC_55_4, I5=>output_MAC_55_5, I6=>output_MAC_55_6, I7=>output_MAC_55_7, I8=>output_MAC_55_8, I9=>output_MAC_55_9, I10=>output_MAC_55_10, I11=>output_MAC_55_11, I12=>output_MAC_55_12, I13=>output_MAC_55_13, I14=>output_MAC_55_14, I15=>output_MAC_55_15, I16=>output_MAC_55_16, I17=>output_MAC_55_17, I18=>output_MAC_55_18, I19=>output_MAC_55_19, I20=>output_MAC_55_20, I21=>output_MAC_55_21, I22=>output_MAC_55_22, I23=>output_MAC_55_23, I24=>output_MAC_55_24, I25=>output_MAC_55_25, I26=>output_MAC_55_26, I27=>output_MAC_55_27, I28=>output_MAC_55_28, I29=>output_MAC_55_29, I30=>output_MAC_55_30, I31=>output_MAC_55_31, 
		SEL_mux=>SEL_mux, O=>output_row_55);

	mux_row_56: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_56_0, I1=>output_MAC_56_1, I2=>output_MAC_56_2, I3=>output_MAC_56_3, I4=>output_MAC_56_4, I5=>output_MAC_56_5, I6=>output_MAC_56_6, I7=>output_MAC_56_7, I8=>output_MAC_56_8, I9=>output_MAC_56_9, I10=>output_MAC_56_10, I11=>output_MAC_56_11, I12=>output_MAC_56_12, I13=>output_MAC_56_13, I14=>output_MAC_56_14, I15=>output_MAC_56_15, I16=>output_MAC_56_16, I17=>output_MAC_56_17, I18=>output_MAC_56_18, I19=>output_MAC_56_19, I20=>output_MAC_56_20, I21=>output_MAC_56_21, I22=>output_MAC_56_22, I23=>output_MAC_56_23, I24=>output_MAC_56_24, I25=>output_MAC_56_25, I26=>output_MAC_56_26, I27=>output_MAC_56_27, I28=>output_MAC_56_28, I29=>output_MAC_56_29, I30=>output_MAC_56_30, I31=>output_MAC_56_31, 
		SEL_mux=>SEL_mux, O=>output_row_56);

	mux_row_57: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_57_0, I1=>output_MAC_57_1, I2=>output_MAC_57_2, I3=>output_MAC_57_3, I4=>output_MAC_57_4, I5=>output_MAC_57_5, I6=>output_MAC_57_6, I7=>output_MAC_57_7, I8=>output_MAC_57_8, I9=>output_MAC_57_9, I10=>output_MAC_57_10, I11=>output_MAC_57_11, I12=>output_MAC_57_12, I13=>output_MAC_57_13, I14=>output_MAC_57_14, I15=>output_MAC_57_15, I16=>output_MAC_57_16, I17=>output_MAC_57_17, I18=>output_MAC_57_18, I19=>output_MAC_57_19, I20=>output_MAC_57_20, I21=>output_MAC_57_21, I22=>output_MAC_57_22, I23=>output_MAC_57_23, I24=>output_MAC_57_24, I25=>output_MAC_57_25, I26=>output_MAC_57_26, I27=>output_MAC_57_27, I28=>output_MAC_57_28, I29=>output_MAC_57_29, I30=>output_MAC_57_30, I31=>output_MAC_57_31, 
		SEL_mux=>SEL_mux, O=>output_row_57);

	mux_row_58: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_58_0, I1=>output_MAC_58_1, I2=>output_MAC_58_2, I3=>output_MAC_58_3, I4=>output_MAC_58_4, I5=>output_MAC_58_5, I6=>output_MAC_58_6, I7=>output_MAC_58_7, I8=>output_MAC_58_8, I9=>output_MAC_58_9, I10=>output_MAC_58_10, I11=>output_MAC_58_11, I12=>output_MAC_58_12, I13=>output_MAC_58_13, I14=>output_MAC_58_14, I15=>output_MAC_58_15, I16=>output_MAC_58_16, I17=>output_MAC_58_17, I18=>output_MAC_58_18, I19=>output_MAC_58_19, I20=>output_MAC_58_20, I21=>output_MAC_58_21, I22=>output_MAC_58_22, I23=>output_MAC_58_23, I24=>output_MAC_58_24, I25=>output_MAC_58_25, I26=>output_MAC_58_26, I27=>output_MAC_58_27, I28=>output_MAC_58_28, I29=>output_MAC_58_29, I30=>output_MAC_58_30, I31=>output_MAC_58_31, 
		SEL_mux=>SEL_mux, O=>output_row_58);

	mux_row_59: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_59_0, I1=>output_MAC_59_1, I2=>output_MAC_59_2, I3=>output_MAC_59_3, I4=>output_MAC_59_4, I5=>output_MAC_59_5, I6=>output_MAC_59_6, I7=>output_MAC_59_7, I8=>output_MAC_59_8, I9=>output_MAC_59_9, I10=>output_MAC_59_10, I11=>output_MAC_59_11, I12=>output_MAC_59_12, I13=>output_MAC_59_13, I14=>output_MAC_59_14, I15=>output_MAC_59_15, I16=>output_MAC_59_16, I17=>output_MAC_59_17, I18=>output_MAC_59_18, I19=>output_MAC_59_19, I20=>output_MAC_59_20, I21=>output_MAC_59_21, I22=>output_MAC_59_22, I23=>output_MAC_59_23, I24=>output_MAC_59_24, I25=>output_MAC_59_25, I26=>output_MAC_59_26, I27=>output_MAC_59_27, I28=>output_MAC_59_28, I29=>output_MAC_59_29, I30=>output_MAC_59_30, I31=>output_MAC_59_31, 
		SEL_mux=>SEL_mux, O=>output_row_59);

	mux_row_60: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_60_0, I1=>output_MAC_60_1, I2=>output_MAC_60_2, I3=>output_MAC_60_3, I4=>output_MAC_60_4, I5=>output_MAC_60_5, I6=>output_MAC_60_6, I7=>output_MAC_60_7, I8=>output_MAC_60_8, I9=>output_MAC_60_9, I10=>output_MAC_60_10, I11=>output_MAC_60_11, I12=>output_MAC_60_12, I13=>output_MAC_60_13, I14=>output_MAC_60_14, I15=>output_MAC_60_15, I16=>output_MAC_60_16, I17=>output_MAC_60_17, I18=>output_MAC_60_18, I19=>output_MAC_60_19, I20=>output_MAC_60_20, I21=>output_MAC_60_21, I22=>output_MAC_60_22, I23=>output_MAC_60_23, I24=>output_MAC_60_24, I25=>output_MAC_60_25, I26=>output_MAC_60_26, I27=>output_MAC_60_27, I28=>output_MAC_60_28, I29=>output_MAC_60_29, I30=>output_MAC_60_30, I31=>output_MAC_60_31, 
		SEL_mux=>SEL_mux, O=>output_row_60);

	mux_row_61: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_61_0, I1=>output_MAC_61_1, I2=>output_MAC_61_2, I3=>output_MAC_61_3, I4=>output_MAC_61_4, I5=>output_MAC_61_5, I6=>output_MAC_61_6, I7=>output_MAC_61_7, I8=>output_MAC_61_8, I9=>output_MAC_61_9, I10=>output_MAC_61_10, I11=>output_MAC_61_11, I12=>output_MAC_61_12, I13=>output_MAC_61_13, I14=>output_MAC_61_14, I15=>output_MAC_61_15, I16=>output_MAC_61_16, I17=>output_MAC_61_17, I18=>output_MAC_61_18, I19=>output_MAC_61_19, I20=>output_MAC_61_20, I21=>output_MAC_61_21, I22=>output_MAC_61_22, I23=>output_MAC_61_23, I24=>output_MAC_61_24, I25=>output_MAC_61_25, I26=>output_MAC_61_26, I27=>output_MAC_61_27, I28=>output_MAC_61_28, I29=>output_MAC_61_29, I30=>output_MAC_61_30, I31=>output_MAC_61_31, 
		SEL_mux=>SEL_mux, O=>output_row_61);

	mux_row_62: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_62_0, I1=>output_MAC_62_1, I2=>output_MAC_62_2, I3=>output_MAC_62_3, I4=>output_MAC_62_4, I5=>output_MAC_62_5, I6=>output_MAC_62_6, I7=>output_MAC_62_7, I8=>output_MAC_62_8, I9=>output_MAC_62_9, I10=>output_MAC_62_10, I11=>output_MAC_62_11, I12=>output_MAC_62_12, I13=>output_MAC_62_13, I14=>output_MAC_62_14, I15=>output_MAC_62_15, I16=>output_MAC_62_16, I17=>output_MAC_62_17, I18=>output_MAC_62_18, I19=>output_MAC_62_19, I20=>output_MAC_62_20, I21=>output_MAC_62_21, I22=>output_MAC_62_22, I23=>output_MAC_62_23, I24=>output_MAC_62_24, I25=>output_MAC_62_25, I26=>output_MAC_62_26, I27=>output_MAC_62_27, I28=>output_MAC_62_28, I29=>output_MAC_62_29, I30=>output_MAC_62_30, I31=>output_MAC_62_31, 
		SEL_mux=>SEL_mux, O=>output_row_62);

	mux_row_63: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_63_0, I1=>output_MAC_63_1, I2=>output_MAC_63_2, I3=>output_MAC_63_3, I4=>output_MAC_63_4, I5=>output_MAC_63_5, I6=>output_MAC_63_6, I7=>output_MAC_63_7, I8=>output_MAC_63_8, I9=>output_MAC_63_9, I10=>output_MAC_63_10, I11=>output_MAC_63_11, I12=>output_MAC_63_12, I13=>output_MAC_63_13, I14=>output_MAC_63_14, I15=>output_MAC_63_15, I16=>output_MAC_63_16, I17=>output_MAC_63_17, I18=>output_MAC_63_18, I19=>output_MAC_63_19, I20=>output_MAC_63_20, I21=>output_MAC_63_21, I22=>output_MAC_63_22, I23=>output_MAC_63_23, I24=>output_MAC_63_24, I25=>output_MAC_63_25, I26=>output_MAC_63_26, I27=>output_MAC_63_27, I28=>output_MAC_63_28, I29=>output_MAC_63_29, I30=>output_MAC_63_30, I31=>output_MAC_63_31, 
		SEL_mux=>SEL_mux, O=>output_row_63);


END behaviour;
