
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MAC_bias_8x768_8 IS
PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7: IN STD_LOGIC_VECTOR(7 downto 0);
	input_col_0, input_col_1, input_col_2, input_col_3, input_col_4, input_col_5, input_col_6, input_col_7, input_col_8, input_col_9, 
	input_col_10, input_col_11, input_col_12, input_col_13, input_col_14, input_col_15, input_col_16, input_col_17, input_col_18, input_col_19, 
	input_col_20, input_col_21, input_col_22, input_col_23, input_col_24, input_col_25, input_col_26, input_col_27, input_col_28, input_col_29, 
	input_col_30, input_col_31, input_col_32, input_col_33, input_col_34, input_col_35, input_col_36, input_col_37, input_col_38, input_col_39, 
	input_col_40, input_col_41, input_col_42, input_col_43, input_col_44, input_col_45, input_col_46, input_col_47, input_col_48, input_col_49, 
	input_col_50, input_col_51, input_col_52, input_col_53, input_col_54, input_col_55, input_col_56, input_col_57, input_col_58, input_col_59, 
	input_col_60, input_col_61, input_col_62, input_col_63, input_col_64, input_col_65, input_col_66, input_col_67, input_col_68, input_col_69, 
	input_col_70, input_col_71, input_col_72, input_col_73, input_col_74, input_col_75, input_col_76, input_col_77, input_col_78, input_col_79, 
	input_col_80, input_col_81, input_col_82, input_col_83, input_col_84, input_col_85, input_col_86, input_col_87, input_col_88, input_col_89, 
	input_col_90, input_col_91, input_col_92, input_col_93, input_col_94, input_col_95, input_col_96, input_col_97, input_col_98, input_col_99, 
	input_col_100, input_col_101, input_col_102, input_col_103, input_col_104, input_col_105, input_col_106, input_col_107, input_col_108, input_col_109, 
	input_col_110, input_col_111, input_col_112, input_col_113, input_col_114, input_col_115, input_col_116, input_col_117, input_col_118, input_col_119, 
	input_col_120, input_col_121, input_col_122, input_col_123, input_col_124, input_col_125, input_col_126, input_col_127, input_col_128, input_col_129, 
	input_col_130, input_col_131, input_col_132, input_col_133, input_col_134, input_col_135, input_col_136, input_col_137, input_col_138, input_col_139, 
	input_col_140, input_col_141, input_col_142, input_col_143, input_col_144, input_col_145, input_col_146, input_col_147, input_col_148, input_col_149, 
	input_col_150, input_col_151, input_col_152, input_col_153, input_col_154, input_col_155, input_col_156, input_col_157, input_col_158, input_col_159, 
	input_col_160, input_col_161, input_col_162, input_col_163, input_col_164, input_col_165, input_col_166, input_col_167, input_col_168, input_col_169, 
	input_col_170, input_col_171, input_col_172, input_col_173, input_col_174, input_col_175, input_col_176, input_col_177, input_col_178, input_col_179, 
	input_col_180, input_col_181, input_col_182, input_col_183, input_col_184, input_col_185, input_col_186, input_col_187, input_col_188, input_col_189, 
	input_col_190, input_col_191, input_col_192, input_col_193, input_col_194, input_col_195, input_col_196, input_col_197, input_col_198, input_col_199, 
	input_col_200, input_col_201, input_col_202, input_col_203, input_col_204, input_col_205, input_col_206, input_col_207, input_col_208, input_col_209, 
	input_col_210, input_col_211, input_col_212, input_col_213, input_col_214, input_col_215, input_col_216, input_col_217, input_col_218, input_col_219, 
	input_col_220, input_col_221, input_col_222, input_col_223, input_col_224, input_col_225, input_col_226, input_col_227, input_col_228, input_col_229, 
	input_col_230, input_col_231, input_col_232, input_col_233, input_col_234, input_col_235, input_col_236, input_col_237, input_col_238, input_col_239, 
	input_col_240, input_col_241, input_col_242, input_col_243, input_col_244, input_col_245, input_col_246, input_col_247, input_col_248, input_col_249, 
	input_col_250, input_col_251, input_col_252, input_col_253, input_col_254, input_col_255, input_col_256, input_col_257, input_col_258, input_col_259, 
	input_col_260, input_col_261, input_col_262, input_col_263, input_col_264, input_col_265, input_col_266, input_col_267, input_col_268, input_col_269, 
	input_col_270, input_col_271, input_col_272, input_col_273, input_col_274, input_col_275, input_col_276, input_col_277, input_col_278, input_col_279, 
	input_col_280, input_col_281, input_col_282, input_col_283, input_col_284, input_col_285, input_col_286, input_col_287, input_col_288, input_col_289, 
	input_col_290, input_col_291, input_col_292, input_col_293, input_col_294, input_col_295, input_col_296, input_col_297, input_col_298, input_col_299, 
	input_col_300, input_col_301, input_col_302, input_col_303, input_col_304, input_col_305, input_col_306, input_col_307, input_col_308, input_col_309, 
	input_col_310, input_col_311, input_col_312, input_col_313, input_col_314, input_col_315, input_col_316, input_col_317, input_col_318, input_col_319, 
	input_col_320, input_col_321, input_col_322, input_col_323, input_col_324, input_col_325, input_col_326, input_col_327, input_col_328, input_col_329, 
	input_col_330, input_col_331, input_col_332, input_col_333, input_col_334, input_col_335, input_col_336, input_col_337, input_col_338, input_col_339, 
	input_col_340, input_col_341, input_col_342, input_col_343, input_col_344, input_col_345, input_col_346, input_col_347, input_col_348, input_col_349, 
	input_col_350, input_col_351, input_col_352, input_col_353, input_col_354, input_col_355, input_col_356, input_col_357, input_col_358, input_col_359, 
	input_col_360, input_col_361, input_col_362, input_col_363, input_col_364, input_col_365, input_col_366, input_col_367, input_col_368, input_col_369, 
	input_col_370, input_col_371, input_col_372, input_col_373, input_col_374, input_col_375, input_col_376, input_col_377, input_col_378, input_col_379, 
	input_col_380, input_col_381, input_col_382, input_col_383, input_col_384, input_col_385, input_col_386, input_col_387, input_col_388, input_col_389, 
	input_col_390, input_col_391, input_col_392, input_col_393, input_col_394, input_col_395, input_col_396, input_col_397, input_col_398, input_col_399, 
	input_col_400, input_col_401, input_col_402, input_col_403, input_col_404, input_col_405, input_col_406, input_col_407, input_col_408, input_col_409, 
	input_col_410, input_col_411, input_col_412, input_col_413, input_col_414, input_col_415, input_col_416, input_col_417, input_col_418, input_col_419, 
	input_col_420, input_col_421, input_col_422, input_col_423, input_col_424, input_col_425, input_col_426, input_col_427, input_col_428, input_col_429, 
	input_col_430, input_col_431, input_col_432, input_col_433, input_col_434, input_col_435, input_col_436, input_col_437, input_col_438, input_col_439, 
	input_col_440, input_col_441, input_col_442, input_col_443, input_col_444, input_col_445, input_col_446, input_col_447, input_col_448, input_col_449, 
	input_col_450, input_col_451, input_col_452, input_col_453, input_col_454, input_col_455, input_col_456, input_col_457, input_col_458, input_col_459, 
	input_col_460, input_col_461, input_col_462, input_col_463, input_col_464, input_col_465, input_col_466, input_col_467, input_col_468, input_col_469, 
	input_col_470, input_col_471, input_col_472, input_col_473, input_col_474, input_col_475, input_col_476, input_col_477, input_col_478, input_col_479, 
	input_col_480, input_col_481, input_col_482, input_col_483, input_col_484, input_col_485, input_col_486, input_col_487, input_col_488, input_col_489, 
	input_col_490, input_col_491, input_col_492, input_col_493, input_col_494, input_col_495, input_col_496, input_col_497, input_col_498, input_col_499, 
	input_col_500, input_col_501, input_col_502, input_col_503, input_col_504, input_col_505, input_col_506, input_col_507, input_col_508, input_col_509, 
	input_col_510, input_col_511, input_col_512, input_col_513, input_col_514, input_col_515, input_col_516, input_col_517, input_col_518, input_col_519, 
	input_col_520, input_col_521, input_col_522, input_col_523, input_col_524, input_col_525, input_col_526, input_col_527, input_col_528, input_col_529, 
	input_col_530, input_col_531, input_col_532, input_col_533, input_col_534, input_col_535, input_col_536, input_col_537, input_col_538, input_col_539, 
	input_col_540, input_col_541, input_col_542, input_col_543, input_col_544, input_col_545, input_col_546, input_col_547, input_col_548, input_col_549, 
	input_col_550, input_col_551, input_col_552, input_col_553, input_col_554, input_col_555, input_col_556, input_col_557, input_col_558, input_col_559, 
	input_col_560, input_col_561, input_col_562, input_col_563, input_col_564, input_col_565, input_col_566, input_col_567, input_col_568, input_col_569, 
	input_col_570, input_col_571, input_col_572, input_col_573, input_col_574, input_col_575, input_col_576, input_col_577, input_col_578, input_col_579, 
	input_col_580, input_col_581, input_col_582, input_col_583, input_col_584, input_col_585, input_col_586, input_col_587, input_col_588, input_col_589, 
	input_col_590, input_col_591, input_col_592, input_col_593, input_col_594, input_col_595, input_col_596, input_col_597, input_col_598, input_col_599, 
	input_col_600, input_col_601, input_col_602, input_col_603, input_col_604, input_col_605, input_col_606, input_col_607, input_col_608, input_col_609, 
	input_col_610, input_col_611, input_col_612, input_col_613, input_col_614, input_col_615, input_col_616, input_col_617, input_col_618, input_col_619, 
	input_col_620, input_col_621, input_col_622, input_col_623, input_col_624, input_col_625, input_col_626, input_col_627, input_col_628, input_col_629, 
	input_col_630, input_col_631, input_col_632, input_col_633, input_col_634, input_col_635, input_col_636, input_col_637, input_col_638, input_col_639, 
	input_col_640, input_col_641, input_col_642, input_col_643, input_col_644, input_col_645, input_col_646, input_col_647, input_col_648, input_col_649, 
	input_col_650, input_col_651, input_col_652, input_col_653, input_col_654, input_col_655, input_col_656, input_col_657, input_col_658, input_col_659, 
	input_col_660, input_col_661, input_col_662, input_col_663, input_col_664, input_col_665, input_col_666, input_col_667, input_col_668, input_col_669, 
	input_col_670, input_col_671, input_col_672, input_col_673, input_col_674, input_col_675, input_col_676, input_col_677, input_col_678, input_col_679, 
	input_col_680, input_col_681, input_col_682, input_col_683, input_col_684, input_col_685, input_col_686, input_col_687, input_col_688, input_col_689, 
	input_col_690, input_col_691, input_col_692, input_col_693, input_col_694, input_col_695, input_col_696, input_col_697, input_col_698, input_col_699, 
	input_col_700, input_col_701, input_col_702, input_col_703, input_col_704, input_col_705, input_col_706, input_col_707, input_col_708, input_col_709, 
	input_col_710, input_col_711, input_col_712, input_col_713, input_col_714, input_col_715, input_col_716, input_col_717, input_col_718, input_col_719, 
	input_col_720, input_col_721, input_col_722, input_col_723, input_col_724, input_col_725, input_col_726, input_col_727, input_col_728, input_col_729, 
	input_col_730, input_col_731, input_col_732, input_col_733, input_col_734, input_col_735, input_col_736, input_col_737, input_col_738, input_col_739, 
	input_col_740, input_col_741, input_col_742, input_col_743, input_col_744, input_col_745, input_col_746, input_col_747, input_col_748, input_col_749, 
	input_col_750, input_col_751, input_col_752, input_col_753, input_col_754, input_col_755, input_col_756, input_col_757, input_col_758, input_col_759, 
	input_col_760, input_col_761, input_col_762, input_col_763, input_col_764, input_col_765, input_col_766, input_col_767: IN STD_LOGIC_VECTOR(7 downto 0);
	b_col : IN STD_LOGIC_VECTOR(31 downto 0);
	SEL_mux: IN STD_LOGIC_VECTOR(9 downto 0);
	CLK, RST_n, ENABLE : IN STD_LOGIC;
	output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7: OUT STD_LOGIC_VECTOR(31 downto 0)
);
END MAC_bias_8x768_8;

ARCHITECTURE behaviour OF  MAC_bias_8x768_8 IS


	COMPONENT MAC_8x768_8 IS
	PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7: IN STD_LOGIC_VECTOR(7 downto 0);
		input_col_0, input_col_1, input_col_2, input_col_3, input_col_4, input_col_5, input_col_6, input_col_7, input_col_8, input_col_9, 
		input_col_10, input_col_11, input_col_12, input_col_13, input_col_14, input_col_15, input_col_16, input_col_17, input_col_18, input_col_19, 
		input_col_20, input_col_21, input_col_22, input_col_23, input_col_24, input_col_25, input_col_26, input_col_27, input_col_28, input_col_29, 
		input_col_30, input_col_31, input_col_32, input_col_33, input_col_34, input_col_35, input_col_36, input_col_37, input_col_38, input_col_39, 
		input_col_40, input_col_41, input_col_42, input_col_43, input_col_44, input_col_45, input_col_46, input_col_47, input_col_48, input_col_49, 
		input_col_50, input_col_51, input_col_52, input_col_53, input_col_54, input_col_55, input_col_56, input_col_57, input_col_58, input_col_59, 
		input_col_60, input_col_61, input_col_62, input_col_63, input_col_64, input_col_65, input_col_66, input_col_67, input_col_68, input_col_69, 
		input_col_70, input_col_71, input_col_72, input_col_73, input_col_74, input_col_75, input_col_76, input_col_77, input_col_78, input_col_79, 
		input_col_80, input_col_81, input_col_82, input_col_83, input_col_84, input_col_85, input_col_86, input_col_87, input_col_88, input_col_89, 
		input_col_90, input_col_91, input_col_92, input_col_93, input_col_94, input_col_95, input_col_96, input_col_97, input_col_98, input_col_99, 
		input_col_100, input_col_101, input_col_102, input_col_103, input_col_104, input_col_105, input_col_106, input_col_107, input_col_108, input_col_109, 
		input_col_110, input_col_111, input_col_112, input_col_113, input_col_114, input_col_115, input_col_116, input_col_117, input_col_118, input_col_119, 
		input_col_120, input_col_121, input_col_122, input_col_123, input_col_124, input_col_125, input_col_126, input_col_127, input_col_128, input_col_129, 
		input_col_130, input_col_131, input_col_132, input_col_133, input_col_134, input_col_135, input_col_136, input_col_137, input_col_138, input_col_139, 
		input_col_140, input_col_141, input_col_142, input_col_143, input_col_144, input_col_145, input_col_146, input_col_147, input_col_148, input_col_149, 
		input_col_150, input_col_151, input_col_152, input_col_153, input_col_154, input_col_155, input_col_156, input_col_157, input_col_158, input_col_159, 
		input_col_160, input_col_161, input_col_162, input_col_163, input_col_164, input_col_165, input_col_166, input_col_167, input_col_168, input_col_169, 
		input_col_170, input_col_171, input_col_172, input_col_173, input_col_174, input_col_175, input_col_176, input_col_177, input_col_178, input_col_179, 
		input_col_180, input_col_181, input_col_182, input_col_183, input_col_184, input_col_185, input_col_186, input_col_187, input_col_188, input_col_189, 
		input_col_190, input_col_191, input_col_192, input_col_193, input_col_194, input_col_195, input_col_196, input_col_197, input_col_198, input_col_199, 
		input_col_200, input_col_201, input_col_202, input_col_203, input_col_204, input_col_205, input_col_206, input_col_207, input_col_208, input_col_209, 
		input_col_210, input_col_211, input_col_212, input_col_213, input_col_214, input_col_215, input_col_216, input_col_217, input_col_218, input_col_219, 
		input_col_220, input_col_221, input_col_222, input_col_223, input_col_224, input_col_225, input_col_226, input_col_227, input_col_228, input_col_229, 
		input_col_230, input_col_231, input_col_232, input_col_233, input_col_234, input_col_235, input_col_236, input_col_237, input_col_238, input_col_239, 
		input_col_240, input_col_241, input_col_242, input_col_243, input_col_244, input_col_245, input_col_246, input_col_247, input_col_248, input_col_249, 
		input_col_250, input_col_251, input_col_252, input_col_253, input_col_254, input_col_255, input_col_256, input_col_257, input_col_258, input_col_259, 
		input_col_260, input_col_261, input_col_262, input_col_263, input_col_264, input_col_265, input_col_266, input_col_267, input_col_268, input_col_269, 
		input_col_270, input_col_271, input_col_272, input_col_273, input_col_274, input_col_275, input_col_276, input_col_277, input_col_278, input_col_279, 
		input_col_280, input_col_281, input_col_282, input_col_283, input_col_284, input_col_285, input_col_286, input_col_287, input_col_288, input_col_289, 
		input_col_290, input_col_291, input_col_292, input_col_293, input_col_294, input_col_295, input_col_296, input_col_297, input_col_298, input_col_299, 
		input_col_300, input_col_301, input_col_302, input_col_303, input_col_304, input_col_305, input_col_306, input_col_307, input_col_308, input_col_309, 
		input_col_310, input_col_311, input_col_312, input_col_313, input_col_314, input_col_315, input_col_316, input_col_317, input_col_318, input_col_319, 
		input_col_320, input_col_321, input_col_322, input_col_323, input_col_324, input_col_325, input_col_326, input_col_327, input_col_328, input_col_329, 
		input_col_330, input_col_331, input_col_332, input_col_333, input_col_334, input_col_335, input_col_336, input_col_337, input_col_338, input_col_339, 
		input_col_340, input_col_341, input_col_342, input_col_343, input_col_344, input_col_345, input_col_346, input_col_347, input_col_348, input_col_349, 
		input_col_350, input_col_351, input_col_352, input_col_353, input_col_354, input_col_355, input_col_356, input_col_357, input_col_358, input_col_359, 
		input_col_360, input_col_361, input_col_362, input_col_363, input_col_364, input_col_365, input_col_366, input_col_367, input_col_368, input_col_369, 
		input_col_370, input_col_371, input_col_372, input_col_373, input_col_374, input_col_375, input_col_376, input_col_377, input_col_378, input_col_379, 
		input_col_380, input_col_381, input_col_382, input_col_383, input_col_384, input_col_385, input_col_386, input_col_387, input_col_388, input_col_389, 
		input_col_390, input_col_391, input_col_392, input_col_393, input_col_394, input_col_395, input_col_396, input_col_397, input_col_398, input_col_399, 
		input_col_400, input_col_401, input_col_402, input_col_403, input_col_404, input_col_405, input_col_406, input_col_407, input_col_408, input_col_409, 
		input_col_410, input_col_411, input_col_412, input_col_413, input_col_414, input_col_415, input_col_416, input_col_417, input_col_418, input_col_419, 
		input_col_420, input_col_421, input_col_422, input_col_423, input_col_424, input_col_425, input_col_426, input_col_427, input_col_428, input_col_429, 
		input_col_430, input_col_431, input_col_432, input_col_433, input_col_434, input_col_435, input_col_436, input_col_437, input_col_438, input_col_439, 
		input_col_440, input_col_441, input_col_442, input_col_443, input_col_444, input_col_445, input_col_446, input_col_447, input_col_448, input_col_449, 
		input_col_450, input_col_451, input_col_452, input_col_453, input_col_454, input_col_455, input_col_456, input_col_457, input_col_458, input_col_459, 
		input_col_460, input_col_461, input_col_462, input_col_463, input_col_464, input_col_465, input_col_466, input_col_467, input_col_468, input_col_469, 
		input_col_470, input_col_471, input_col_472, input_col_473, input_col_474, input_col_475, input_col_476, input_col_477, input_col_478, input_col_479, 
		input_col_480, input_col_481, input_col_482, input_col_483, input_col_484, input_col_485, input_col_486, input_col_487, input_col_488, input_col_489, 
		input_col_490, input_col_491, input_col_492, input_col_493, input_col_494, input_col_495, input_col_496, input_col_497, input_col_498, input_col_499, 
		input_col_500, input_col_501, input_col_502, input_col_503, input_col_504, input_col_505, input_col_506, input_col_507, input_col_508, input_col_509, 
		input_col_510, input_col_511, input_col_512, input_col_513, input_col_514, input_col_515, input_col_516, input_col_517, input_col_518, input_col_519, 
		input_col_520, input_col_521, input_col_522, input_col_523, input_col_524, input_col_525, input_col_526, input_col_527, input_col_528, input_col_529, 
		input_col_530, input_col_531, input_col_532, input_col_533, input_col_534, input_col_535, input_col_536, input_col_537, input_col_538, input_col_539, 
		input_col_540, input_col_541, input_col_542, input_col_543, input_col_544, input_col_545, input_col_546, input_col_547, input_col_548, input_col_549, 
		input_col_550, input_col_551, input_col_552, input_col_553, input_col_554, input_col_555, input_col_556, input_col_557, input_col_558, input_col_559, 
		input_col_560, input_col_561, input_col_562, input_col_563, input_col_564, input_col_565, input_col_566, input_col_567, input_col_568, input_col_569, 
		input_col_570, input_col_571, input_col_572, input_col_573, input_col_574, input_col_575, input_col_576, input_col_577, input_col_578, input_col_579, 
		input_col_580, input_col_581, input_col_582, input_col_583, input_col_584, input_col_585, input_col_586, input_col_587, input_col_588, input_col_589, 
		input_col_590, input_col_591, input_col_592, input_col_593, input_col_594, input_col_595, input_col_596, input_col_597, input_col_598, input_col_599, 
		input_col_600, input_col_601, input_col_602, input_col_603, input_col_604, input_col_605, input_col_606, input_col_607, input_col_608, input_col_609, 
		input_col_610, input_col_611, input_col_612, input_col_613, input_col_614, input_col_615, input_col_616, input_col_617, input_col_618, input_col_619, 
		input_col_620, input_col_621, input_col_622, input_col_623, input_col_624, input_col_625, input_col_626, input_col_627, input_col_628, input_col_629, 
		input_col_630, input_col_631, input_col_632, input_col_633, input_col_634, input_col_635, input_col_636, input_col_637, input_col_638, input_col_639, 
		input_col_640, input_col_641, input_col_642, input_col_643, input_col_644, input_col_645, input_col_646, input_col_647, input_col_648, input_col_649, 
		input_col_650, input_col_651, input_col_652, input_col_653, input_col_654, input_col_655, input_col_656, input_col_657, input_col_658, input_col_659, 
		input_col_660, input_col_661, input_col_662, input_col_663, input_col_664, input_col_665, input_col_666, input_col_667, input_col_668, input_col_669, 
		input_col_670, input_col_671, input_col_672, input_col_673, input_col_674, input_col_675, input_col_676, input_col_677, input_col_678, input_col_679, 
		input_col_680, input_col_681, input_col_682, input_col_683, input_col_684, input_col_685, input_col_686, input_col_687, input_col_688, input_col_689, 
		input_col_690, input_col_691, input_col_692, input_col_693, input_col_694, input_col_695, input_col_696, input_col_697, input_col_698, input_col_699, 
		input_col_700, input_col_701, input_col_702, input_col_703, input_col_704, input_col_705, input_col_706, input_col_707, input_col_708, input_col_709, 
		input_col_710, input_col_711, input_col_712, input_col_713, input_col_714, input_col_715, input_col_716, input_col_717, input_col_718, input_col_719, 
		input_col_720, input_col_721, input_col_722, input_col_723, input_col_724, input_col_725, input_col_726, input_col_727, input_col_728, input_col_729, 
		input_col_730, input_col_731, input_col_732, input_col_733, input_col_734, input_col_735, input_col_736, input_col_737, input_col_738, input_col_739, 
		input_col_740, input_col_741, input_col_742, input_col_743, input_col_744, input_col_745, input_col_746, input_col_747, input_col_748, input_col_749, 
		input_col_750, input_col_751, input_col_752, input_col_753, input_col_754, input_col_755, input_col_756, input_col_757, input_col_758, input_col_759, 
		input_col_760, input_col_761, input_col_762, input_col_763, input_col_764, input_col_765, input_col_766, input_col_767: IN STD_LOGIC_VECTOR(7 downto 0);
		SEL_mux: IN STD_LOGIC_VECTOR(9 downto 0);
		CLK, RST_n, ENABLE : IN STD_LOGIC;
		output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7: OUT STD_LOGIC_VECTOR(31 downto 0)
	);
	END COMPONENT;


	COMPONENT bias_sum_8_32 IS
	PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7: IN STD_LOGIC_VECTOR(31 downto 0);
		b_col : IN STD_LOGIC_VECTOR(31 downto 0);
		output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7: OUT STD_LOGIC_VECTOR(31 downto 0)
	);
	END COMPONENT;


	SIGNAL output_row_MAC_base_0: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_row_MAC_base_1: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_row_MAC_base_2: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_row_MAC_base_3: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_row_MAC_base_4: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_row_MAC_base_5: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_row_MAC_base_6: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_row_MAC_base_7: STD_LOGIC_VECTOR(31 downto 0);

BEGIN

	MAC_base: MAC_8x768_8 PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE,
		input_row_0=>input_row_0, input_row_1=>input_row_1, input_row_2=>input_row_2, input_row_3=>input_row_3, input_row_4=>input_row_4, input_row_5=>input_row_5, input_row_6=>input_row_6, input_row_7=>input_row_7, 
		input_col_0=>input_col_0, input_col_1=>input_col_1, input_col_2=>input_col_2, input_col_3=>input_col_3, input_col_4=>input_col_4, input_col_5=>input_col_5, input_col_6=>input_col_6, input_col_7=>input_col_7, input_col_8=>input_col_8, input_col_9=>input_col_9, input_col_10=>input_col_10, input_col_11=>input_col_11, input_col_12=>input_col_12, input_col_13=>input_col_13, input_col_14=>input_col_14, input_col_15=>input_col_15, input_col_16=>input_col_16, input_col_17=>input_col_17, input_col_18=>input_col_18, input_col_19=>input_col_19, input_col_20=>input_col_20, input_col_21=>input_col_21, input_col_22=>input_col_22, input_col_23=>input_col_23, input_col_24=>input_col_24, input_col_25=>input_col_25, input_col_26=>input_col_26, input_col_27=>input_col_27, input_col_28=>input_col_28, input_col_29=>input_col_29, input_col_30=>input_col_30, input_col_31=>input_col_31, input_col_32=>input_col_32, input_col_33=>input_col_33, input_col_34=>input_col_34, input_col_35=>input_col_35, input_col_36=>input_col_36, input_col_37=>input_col_37, input_col_38=>input_col_38, input_col_39=>input_col_39, input_col_40=>input_col_40, input_col_41=>input_col_41, input_col_42=>input_col_42, input_col_43=>input_col_43, input_col_44=>input_col_44, input_col_45=>input_col_45, input_col_46=>input_col_46, input_col_47=>input_col_47, input_col_48=>input_col_48, input_col_49=>input_col_49, input_col_50=>input_col_50, input_col_51=>input_col_51, input_col_52=>input_col_52, input_col_53=>input_col_53, input_col_54=>input_col_54, input_col_55=>input_col_55, input_col_56=>input_col_56, input_col_57=>input_col_57, input_col_58=>input_col_58, input_col_59=>input_col_59, input_col_60=>input_col_60, input_col_61=>input_col_61, input_col_62=>input_col_62, input_col_63=>input_col_63, input_col_64=>input_col_64, input_col_65=>input_col_65, input_col_66=>input_col_66, input_col_67=>input_col_67, input_col_68=>input_col_68, input_col_69=>input_col_69, input_col_70=>input_col_70, input_col_71=>input_col_71, input_col_72=>input_col_72, input_col_73=>input_col_73, input_col_74=>input_col_74, input_col_75=>input_col_75, input_col_76=>input_col_76, input_col_77=>input_col_77, input_col_78=>input_col_78, input_col_79=>input_col_79, input_col_80=>input_col_80, input_col_81=>input_col_81, input_col_82=>input_col_82, input_col_83=>input_col_83, input_col_84=>input_col_84, input_col_85=>input_col_85, input_col_86=>input_col_86, input_col_87=>input_col_87, input_col_88=>input_col_88, input_col_89=>input_col_89, input_col_90=>input_col_90, input_col_91=>input_col_91, input_col_92=>input_col_92, input_col_93=>input_col_93, input_col_94=>input_col_94, input_col_95=>input_col_95, input_col_96=>input_col_96, input_col_97=>input_col_97, input_col_98=>input_col_98, input_col_99=>input_col_99, input_col_100=>input_col_100, input_col_101=>input_col_101, input_col_102=>input_col_102, input_col_103=>input_col_103, input_col_104=>input_col_104, input_col_105=>input_col_105, input_col_106=>input_col_106, input_col_107=>input_col_107, input_col_108=>input_col_108, input_col_109=>input_col_109, input_col_110=>input_col_110, input_col_111=>input_col_111, input_col_112=>input_col_112, input_col_113=>input_col_113, input_col_114=>input_col_114, input_col_115=>input_col_115, input_col_116=>input_col_116, input_col_117=>input_col_117, input_col_118=>input_col_118, input_col_119=>input_col_119, input_col_120=>input_col_120, input_col_121=>input_col_121, input_col_122=>input_col_122, input_col_123=>input_col_123, input_col_124=>input_col_124, input_col_125=>input_col_125, input_col_126=>input_col_126, input_col_127=>input_col_127, input_col_128=>input_col_128, input_col_129=>input_col_129, input_col_130=>input_col_130, input_col_131=>input_col_131, input_col_132=>input_col_132, input_col_133=>input_col_133, input_col_134=>input_col_134, input_col_135=>input_col_135, input_col_136=>input_col_136, input_col_137=>input_col_137, input_col_138=>input_col_138, input_col_139=>input_col_139, input_col_140=>input_col_140, input_col_141=>input_col_141, input_col_142=>input_col_142, input_col_143=>input_col_143, input_col_144=>input_col_144, input_col_145=>input_col_145, input_col_146=>input_col_146, input_col_147=>input_col_147, input_col_148=>input_col_148, input_col_149=>input_col_149, input_col_150=>input_col_150, input_col_151=>input_col_151, input_col_152=>input_col_152, input_col_153=>input_col_153, input_col_154=>input_col_154, input_col_155=>input_col_155, input_col_156=>input_col_156, input_col_157=>input_col_157, input_col_158=>input_col_158, input_col_159=>input_col_159, input_col_160=>input_col_160, input_col_161=>input_col_161, input_col_162=>input_col_162, input_col_163=>input_col_163, input_col_164=>input_col_164, input_col_165=>input_col_165, input_col_166=>input_col_166, input_col_167=>input_col_167, input_col_168=>input_col_168, input_col_169=>input_col_169, input_col_170=>input_col_170, input_col_171=>input_col_171, input_col_172=>input_col_172, input_col_173=>input_col_173, input_col_174=>input_col_174, input_col_175=>input_col_175, input_col_176=>input_col_176, input_col_177=>input_col_177, input_col_178=>input_col_178, input_col_179=>input_col_179, input_col_180=>input_col_180, input_col_181=>input_col_181, input_col_182=>input_col_182, input_col_183=>input_col_183, input_col_184=>input_col_184, input_col_185=>input_col_185, input_col_186=>input_col_186, input_col_187=>input_col_187, input_col_188=>input_col_188, input_col_189=>input_col_189, input_col_190=>input_col_190, input_col_191=>input_col_191, input_col_192=>input_col_192, input_col_193=>input_col_193, input_col_194=>input_col_194, input_col_195=>input_col_195, input_col_196=>input_col_196, input_col_197=>input_col_197, input_col_198=>input_col_198, input_col_199=>input_col_199, input_col_200=>input_col_200, input_col_201=>input_col_201, input_col_202=>input_col_202, input_col_203=>input_col_203, input_col_204=>input_col_204, input_col_205=>input_col_205, input_col_206=>input_col_206, input_col_207=>input_col_207, input_col_208=>input_col_208, input_col_209=>input_col_209, input_col_210=>input_col_210, input_col_211=>input_col_211, input_col_212=>input_col_212, input_col_213=>input_col_213, input_col_214=>input_col_214, input_col_215=>input_col_215, input_col_216=>input_col_216, input_col_217=>input_col_217, input_col_218=>input_col_218, input_col_219=>input_col_219, input_col_220=>input_col_220, input_col_221=>input_col_221, input_col_222=>input_col_222, input_col_223=>input_col_223, input_col_224=>input_col_224, input_col_225=>input_col_225, input_col_226=>input_col_226, input_col_227=>input_col_227, input_col_228=>input_col_228, input_col_229=>input_col_229, input_col_230=>input_col_230, input_col_231=>input_col_231, input_col_232=>input_col_232, input_col_233=>input_col_233, input_col_234=>input_col_234, input_col_235=>input_col_235, input_col_236=>input_col_236, input_col_237=>input_col_237, input_col_238=>input_col_238, input_col_239=>input_col_239, input_col_240=>input_col_240, input_col_241=>input_col_241, input_col_242=>input_col_242, input_col_243=>input_col_243, input_col_244=>input_col_244, input_col_245=>input_col_245, input_col_246=>input_col_246, input_col_247=>input_col_247, input_col_248=>input_col_248, input_col_249=>input_col_249, input_col_250=>input_col_250, input_col_251=>input_col_251, input_col_252=>input_col_252, input_col_253=>input_col_253, input_col_254=>input_col_254, input_col_255=>input_col_255, input_col_256=>input_col_256, input_col_257=>input_col_257, input_col_258=>input_col_258, input_col_259=>input_col_259, input_col_260=>input_col_260, input_col_261=>input_col_261, input_col_262=>input_col_262, input_col_263=>input_col_263, input_col_264=>input_col_264, input_col_265=>input_col_265, input_col_266=>input_col_266, input_col_267=>input_col_267, input_col_268=>input_col_268, input_col_269=>input_col_269, input_col_270=>input_col_270, input_col_271=>input_col_271, input_col_272=>input_col_272, input_col_273=>input_col_273, input_col_274=>input_col_274, input_col_275=>input_col_275, input_col_276=>input_col_276, input_col_277=>input_col_277, input_col_278=>input_col_278, input_col_279=>input_col_279, input_col_280=>input_col_280, input_col_281=>input_col_281, input_col_282=>input_col_282, input_col_283=>input_col_283, input_col_284=>input_col_284, input_col_285=>input_col_285, input_col_286=>input_col_286, input_col_287=>input_col_287, input_col_288=>input_col_288, input_col_289=>input_col_289, input_col_290=>input_col_290, input_col_291=>input_col_291, input_col_292=>input_col_292, input_col_293=>input_col_293, input_col_294=>input_col_294, input_col_295=>input_col_295, input_col_296=>input_col_296, input_col_297=>input_col_297, input_col_298=>input_col_298, input_col_299=>input_col_299, input_col_300=>input_col_300, input_col_301=>input_col_301, input_col_302=>input_col_302, input_col_303=>input_col_303, input_col_304=>input_col_304, input_col_305=>input_col_305, input_col_306=>input_col_306, input_col_307=>input_col_307, input_col_308=>input_col_308, input_col_309=>input_col_309, input_col_310=>input_col_310, input_col_311=>input_col_311, input_col_312=>input_col_312, input_col_313=>input_col_313, input_col_314=>input_col_314, input_col_315=>input_col_315, input_col_316=>input_col_316, input_col_317=>input_col_317, input_col_318=>input_col_318, input_col_319=>input_col_319, input_col_320=>input_col_320, input_col_321=>input_col_321, input_col_322=>input_col_322, input_col_323=>input_col_323, input_col_324=>input_col_324, input_col_325=>input_col_325, input_col_326=>input_col_326, input_col_327=>input_col_327, input_col_328=>input_col_328, input_col_329=>input_col_329, input_col_330=>input_col_330, input_col_331=>input_col_331, input_col_332=>input_col_332, input_col_333=>input_col_333, input_col_334=>input_col_334, input_col_335=>input_col_335, input_col_336=>input_col_336, input_col_337=>input_col_337, input_col_338=>input_col_338, input_col_339=>input_col_339, input_col_340=>input_col_340, input_col_341=>input_col_341, input_col_342=>input_col_342, input_col_343=>input_col_343, input_col_344=>input_col_344, input_col_345=>input_col_345, input_col_346=>input_col_346, input_col_347=>input_col_347, input_col_348=>input_col_348, input_col_349=>input_col_349, input_col_350=>input_col_350, input_col_351=>input_col_351, input_col_352=>input_col_352, input_col_353=>input_col_353, input_col_354=>input_col_354, input_col_355=>input_col_355, input_col_356=>input_col_356, input_col_357=>input_col_357, input_col_358=>input_col_358, input_col_359=>input_col_359, input_col_360=>input_col_360, input_col_361=>input_col_361, input_col_362=>input_col_362, input_col_363=>input_col_363, input_col_364=>input_col_364, input_col_365=>input_col_365, input_col_366=>input_col_366, input_col_367=>input_col_367, input_col_368=>input_col_368, input_col_369=>input_col_369, input_col_370=>input_col_370, input_col_371=>input_col_371, input_col_372=>input_col_372, input_col_373=>input_col_373, input_col_374=>input_col_374, input_col_375=>input_col_375, input_col_376=>input_col_376, input_col_377=>input_col_377, input_col_378=>input_col_378, input_col_379=>input_col_379, input_col_380=>input_col_380, input_col_381=>input_col_381, input_col_382=>input_col_382, input_col_383=>input_col_383, input_col_384=>input_col_384, input_col_385=>input_col_385, input_col_386=>input_col_386, input_col_387=>input_col_387, input_col_388=>input_col_388, input_col_389=>input_col_389, input_col_390=>input_col_390, input_col_391=>input_col_391, input_col_392=>input_col_392, input_col_393=>input_col_393, input_col_394=>input_col_394, input_col_395=>input_col_395, input_col_396=>input_col_396, input_col_397=>input_col_397, input_col_398=>input_col_398, input_col_399=>input_col_399, input_col_400=>input_col_400, input_col_401=>input_col_401, input_col_402=>input_col_402, input_col_403=>input_col_403, input_col_404=>input_col_404, input_col_405=>input_col_405, input_col_406=>input_col_406, input_col_407=>input_col_407, input_col_408=>input_col_408, input_col_409=>input_col_409, input_col_410=>input_col_410, input_col_411=>input_col_411, input_col_412=>input_col_412, input_col_413=>input_col_413, input_col_414=>input_col_414, input_col_415=>input_col_415, input_col_416=>input_col_416, input_col_417=>input_col_417, input_col_418=>input_col_418, input_col_419=>input_col_419, input_col_420=>input_col_420, input_col_421=>input_col_421, input_col_422=>input_col_422, input_col_423=>input_col_423, input_col_424=>input_col_424, input_col_425=>input_col_425, input_col_426=>input_col_426, input_col_427=>input_col_427, input_col_428=>input_col_428, input_col_429=>input_col_429, input_col_430=>input_col_430, input_col_431=>input_col_431, input_col_432=>input_col_432, input_col_433=>input_col_433, input_col_434=>input_col_434, input_col_435=>input_col_435, input_col_436=>input_col_436, input_col_437=>input_col_437, input_col_438=>input_col_438, input_col_439=>input_col_439, input_col_440=>input_col_440, input_col_441=>input_col_441, input_col_442=>input_col_442, input_col_443=>input_col_443, input_col_444=>input_col_444, input_col_445=>input_col_445, input_col_446=>input_col_446, input_col_447=>input_col_447, input_col_448=>input_col_448, input_col_449=>input_col_449, input_col_450=>input_col_450, input_col_451=>input_col_451, input_col_452=>input_col_452, input_col_453=>input_col_453, input_col_454=>input_col_454, input_col_455=>input_col_455, input_col_456=>input_col_456, input_col_457=>input_col_457, input_col_458=>input_col_458, input_col_459=>input_col_459, input_col_460=>input_col_460, input_col_461=>input_col_461, input_col_462=>input_col_462, input_col_463=>input_col_463, input_col_464=>input_col_464, input_col_465=>input_col_465, input_col_466=>input_col_466, input_col_467=>input_col_467, input_col_468=>input_col_468, input_col_469=>input_col_469, input_col_470=>input_col_470, input_col_471=>input_col_471, input_col_472=>input_col_472, input_col_473=>input_col_473, input_col_474=>input_col_474, input_col_475=>input_col_475, input_col_476=>input_col_476, input_col_477=>input_col_477, input_col_478=>input_col_478, input_col_479=>input_col_479, input_col_480=>input_col_480, input_col_481=>input_col_481, input_col_482=>input_col_482, input_col_483=>input_col_483, input_col_484=>input_col_484, input_col_485=>input_col_485, input_col_486=>input_col_486, input_col_487=>input_col_487, input_col_488=>input_col_488, input_col_489=>input_col_489, input_col_490=>input_col_490, input_col_491=>input_col_491, input_col_492=>input_col_492, input_col_493=>input_col_493, input_col_494=>input_col_494, input_col_495=>input_col_495, input_col_496=>input_col_496, input_col_497=>input_col_497, input_col_498=>input_col_498, input_col_499=>input_col_499, input_col_500=>input_col_500, input_col_501=>input_col_501, input_col_502=>input_col_502, input_col_503=>input_col_503, input_col_504=>input_col_504, input_col_505=>input_col_505, input_col_506=>input_col_506, input_col_507=>input_col_507, input_col_508=>input_col_508, input_col_509=>input_col_509, input_col_510=>input_col_510, input_col_511=>input_col_511, input_col_512=>input_col_512, input_col_513=>input_col_513, input_col_514=>input_col_514, input_col_515=>input_col_515, input_col_516=>input_col_516, input_col_517=>input_col_517, input_col_518=>input_col_518, input_col_519=>input_col_519, input_col_520=>input_col_520, input_col_521=>input_col_521, input_col_522=>input_col_522, input_col_523=>input_col_523, input_col_524=>input_col_524, input_col_525=>input_col_525, input_col_526=>input_col_526, input_col_527=>input_col_527, input_col_528=>input_col_528, input_col_529=>input_col_529, input_col_530=>input_col_530, input_col_531=>input_col_531, input_col_532=>input_col_532, input_col_533=>input_col_533, input_col_534=>input_col_534, input_col_535=>input_col_535, input_col_536=>input_col_536, input_col_537=>input_col_537, input_col_538=>input_col_538, input_col_539=>input_col_539, input_col_540=>input_col_540, input_col_541=>input_col_541, input_col_542=>input_col_542, input_col_543=>input_col_543, input_col_544=>input_col_544, input_col_545=>input_col_545, input_col_546=>input_col_546, input_col_547=>input_col_547, input_col_548=>input_col_548, input_col_549=>input_col_549, input_col_550=>input_col_550, input_col_551=>input_col_551, input_col_552=>input_col_552, input_col_553=>input_col_553, input_col_554=>input_col_554, input_col_555=>input_col_555, input_col_556=>input_col_556, input_col_557=>input_col_557, input_col_558=>input_col_558, input_col_559=>input_col_559, input_col_560=>input_col_560, input_col_561=>input_col_561, input_col_562=>input_col_562, input_col_563=>input_col_563, input_col_564=>input_col_564, input_col_565=>input_col_565, input_col_566=>input_col_566, input_col_567=>input_col_567, input_col_568=>input_col_568, input_col_569=>input_col_569, input_col_570=>input_col_570, input_col_571=>input_col_571, input_col_572=>input_col_572, input_col_573=>input_col_573, input_col_574=>input_col_574, input_col_575=>input_col_575, input_col_576=>input_col_576, input_col_577=>input_col_577, input_col_578=>input_col_578, input_col_579=>input_col_579, input_col_580=>input_col_580, input_col_581=>input_col_581, input_col_582=>input_col_582, input_col_583=>input_col_583, input_col_584=>input_col_584, input_col_585=>input_col_585, input_col_586=>input_col_586, input_col_587=>input_col_587, input_col_588=>input_col_588, input_col_589=>input_col_589, input_col_590=>input_col_590, input_col_591=>input_col_591, input_col_592=>input_col_592, input_col_593=>input_col_593, input_col_594=>input_col_594, input_col_595=>input_col_595, input_col_596=>input_col_596, input_col_597=>input_col_597, input_col_598=>input_col_598, input_col_599=>input_col_599, input_col_600=>input_col_600, input_col_601=>input_col_601, input_col_602=>input_col_602, input_col_603=>input_col_603, input_col_604=>input_col_604, input_col_605=>input_col_605, input_col_606=>input_col_606, input_col_607=>input_col_607, input_col_608=>input_col_608, input_col_609=>input_col_609, input_col_610=>input_col_610, input_col_611=>input_col_611, input_col_612=>input_col_612, input_col_613=>input_col_613, input_col_614=>input_col_614, input_col_615=>input_col_615, input_col_616=>input_col_616, input_col_617=>input_col_617, input_col_618=>input_col_618, input_col_619=>input_col_619, input_col_620=>input_col_620, input_col_621=>input_col_621, input_col_622=>input_col_622, input_col_623=>input_col_623, input_col_624=>input_col_624, input_col_625=>input_col_625, input_col_626=>input_col_626, input_col_627=>input_col_627, input_col_628=>input_col_628, input_col_629=>input_col_629, input_col_630=>input_col_630, input_col_631=>input_col_631, input_col_632=>input_col_632, input_col_633=>input_col_633, input_col_634=>input_col_634, input_col_635=>input_col_635, input_col_636=>input_col_636, input_col_637=>input_col_637, input_col_638=>input_col_638, input_col_639=>input_col_639, input_col_640=>input_col_640, input_col_641=>input_col_641, input_col_642=>input_col_642, input_col_643=>input_col_643, input_col_644=>input_col_644, input_col_645=>input_col_645, input_col_646=>input_col_646, input_col_647=>input_col_647, input_col_648=>input_col_648, input_col_649=>input_col_649, input_col_650=>input_col_650, input_col_651=>input_col_651, input_col_652=>input_col_652, input_col_653=>input_col_653, input_col_654=>input_col_654, input_col_655=>input_col_655, input_col_656=>input_col_656, input_col_657=>input_col_657, input_col_658=>input_col_658, input_col_659=>input_col_659, input_col_660=>input_col_660, input_col_661=>input_col_661, input_col_662=>input_col_662, input_col_663=>input_col_663, input_col_664=>input_col_664, input_col_665=>input_col_665, input_col_666=>input_col_666, input_col_667=>input_col_667, input_col_668=>input_col_668, input_col_669=>input_col_669, input_col_670=>input_col_670, input_col_671=>input_col_671, input_col_672=>input_col_672, input_col_673=>input_col_673, input_col_674=>input_col_674, input_col_675=>input_col_675, input_col_676=>input_col_676, input_col_677=>input_col_677, input_col_678=>input_col_678, input_col_679=>input_col_679, input_col_680=>input_col_680, input_col_681=>input_col_681, input_col_682=>input_col_682, input_col_683=>input_col_683, input_col_684=>input_col_684, input_col_685=>input_col_685, input_col_686=>input_col_686, input_col_687=>input_col_687, input_col_688=>input_col_688, input_col_689=>input_col_689, input_col_690=>input_col_690, input_col_691=>input_col_691, input_col_692=>input_col_692, input_col_693=>input_col_693, input_col_694=>input_col_694, input_col_695=>input_col_695, input_col_696=>input_col_696, input_col_697=>input_col_697, input_col_698=>input_col_698, input_col_699=>input_col_699, input_col_700=>input_col_700, input_col_701=>input_col_701, input_col_702=>input_col_702, input_col_703=>input_col_703, input_col_704=>input_col_704, input_col_705=>input_col_705, input_col_706=>input_col_706, input_col_707=>input_col_707, input_col_708=>input_col_708, input_col_709=>input_col_709, input_col_710=>input_col_710, input_col_711=>input_col_711, input_col_712=>input_col_712, input_col_713=>input_col_713, input_col_714=>input_col_714, input_col_715=>input_col_715, input_col_716=>input_col_716, input_col_717=>input_col_717, input_col_718=>input_col_718, input_col_719=>input_col_719, input_col_720=>input_col_720, input_col_721=>input_col_721, input_col_722=>input_col_722, input_col_723=>input_col_723, input_col_724=>input_col_724, input_col_725=>input_col_725, input_col_726=>input_col_726, input_col_727=>input_col_727, input_col_728=>input_col_728, input_col_729=>input_col_729, input_col_730=>input_col_730, input_col_731=>input_col_731, input_col_732=>input_col_732, input_col_733=>input_col_733, input_col_734=>input_col_734, input_col_735=>input_col_735, input_col_736=>input_col_736, input_col_737=>input_col_737, input_col_738=>input_col_738, input_col_739=>input_col_739, input_col_740=>input_col_740, input_col_741=>input_col_741, input_col_742=>input_col_742, input_col_743=>input_col_743, input_col_744=>input_col_744, input_col_745=>input_col_745, input_col_746=>input_col_746, input_col_747=>input_col_747, input_col_748=>input_col_748, input_col_749=>input_col_749, input_col_750=>input_col_750, input_col_751=>input_col_751, input_col_752=>input_col_752, input_col_753=>input_col_753, input_col_754=>input_col_754, input_col_755=>input_col_755, input_col_756=>input_col_756, input_col_757=>input_col_757, input_col_758=>input_col_758, input_col_759=>input_col_759, input_col_760=>input_col_760, input_col_761=>input_col_761, input_col_762=>input_col_762, input_col_763=>input_col_763, input_col_764=>input_col_764, input_col_765=>input_col_765, input_col_766=>input_col_766, input_col_767=>input_col_767, 
		output_row_0=>output_row_MAC_base_0, output_row_1=>output_row_MAC_base_1, output_row_2=>output_row_MAC_base_2, output_row_3=>output_row_MAC_base_3, output_row_4=>output_row_MAC_base_4, output_row_5=>output_row_MAC_base_5, output_row_6=>output_row_MAC_base_6, output_row_7=>output_row_MAC_base_7, 
		SEL_mux=>SEL_mux);
	bias_sum: bias_sum_8_32 PORT MAP(input_row_0=>output_row_MAC_base_0, input_row_1=>output_row_MAC_base_1, input_row_2=>output_row_MAC_base_2, input_row_3=>output_row_MAC_base_3, input_row_4=>output_row_MAC_base_4, input_row_5=>output_row_MAC_base_5, input_row_6=>output_row_MAC_base_6, input_row_7=>output_row_MAC_base_7, 
		b_col=>b_col, output_row_0=>output_row_0, output_row_1=>output_row_1, output_row_2=>output_row_2, output_row_3=>output_row_3, output_row_4=>output_row_4, output_row_5=>output_row_5, output_row_6=>output_row_6, output_row_7=>output_row_7);


END behaviour;
