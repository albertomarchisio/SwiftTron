
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MAC_64x16_8 IS
PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7, input_row_8, input_row_9, 
	input_row_10, input_row_11, input_row_12, input_row_13, input_row_14, input_row_15, input_row_16, input_row_17, input_row_18, input_row_19, 
	input_row_20, input_row_21, input_row_22, input_row_23, input_row_24, input_row_25, input_row_26, input_row_27, input_row_28, input_row_29, 
	input_row_30, input_row_31, input_row_32, input_row_33, input_row_34, input_row_35, input_row_36, input_row_37, input_row_38, input_row_39, 
	input_row_40, input_row_41, input_row_42, input_row_43, input_row_44, input_row_45, input_row_46, input_row_47, input_row_48, input_row_49, 
	input_row_50, input_row_51, input_row_52, input_row_53, input_row_54, input_row_55, input_row_56, input_row_57, input_row_58, input_row_59, 
	input_row_60, input_row_61, input_row_62, input_row_63: IN STD_LOGIC_VECTOR(7 downto 0);
	input_col_0, input_col_1, input_col_2, input_col_3, input_col_4, input_col_5, input_col_6, input_col_7, input_col_8, input_col_9, 
	input_col_10, input_col_11, input_col_12, input_col_13, input_col_14, input_col_15: IN STD_LOGIC_VECTOR(7 downto 0);
	SEL_mux: IN STD_LOGIC_VECTOR(3 downto 0);
	CLK, RST_n, ENABLE : IN STD_LOGIC;
	output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7, output_row_8, output_row_9, 
	output_row_10, output_row_11, output_row_12, output_row_13, output_row_14, output_row_15, output_row_16, output_row_17, output_row_18, output_row_19, 
	output_row_20, output_row_21, output_row_22, output_row_23, output_row_24, output_row_25, output_row_26, output_row_27, output_row_28, output_row_29, 
	output_row_30, output_row_31, output_row_32, output_row_33, output_row_34, output_row_35, output_row_36, output_row_37, output_row_38, output_row_39, 
	output_row_40, output_row_41, output_row_42, output_row_43, output_row_44, output_row_45, output_row_46, output_row_47, output_row_48, output_row_49, 
	output_row_50, output_row_51, output_row_52, output_row_53, output_row_54, output_row_55, output_row_56, output_row_57, output_row_58, output_row_59, 
	output_row_60, output_row_61, output_row_62, output_row_63: OUT STD_LOGIC_VECTOR(31 downto 0)
);
END MAC_64x16_8;

ARCHITECTURE behaviour OF  MAC_64x16_8 IS

	COMPONENT MAC IS
	GENERIC (data_size : POSITIVE := 2;
	 acc_size : POSITIVE := 16 );
	PORT( data_in_A, data_in_B  : IN STD_LOGIC_VECTOR(data_size-1 downto 0);
		CLK, RST_n, ENABLE 	: IN STD_LOGIC;
		data_out    			: OUT STD_LOGIC_VECTOR(acc_size-1 downto 0));
	END COMPONENT;

	COMPONENT mux_16to1_nbit IS
	GENERIC ( N : POSITIVE :=2);
	PORT(
		I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, 
		I10, I11, I12, I13, I14, I15: IN STD_LOGIC_VECTOR(N-1 downto 0);
		SEL_mux  : IN STD_LOGIC_VECTOR(3 downto 0);
		O    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
	END COMPONENT;


	SIGNAL output_MAC_0_0, output_MAC_0_1, output_MAC_0_2, output_MAC_0_3, output_MAC_0_4, output_MAC_0_5, output_MAC_0_6, output_MAC_0_7, output_MAC_0_8, output_MAC_0_9, 
		output_MAC_0_10, output_MAC_0_11, output_MAC_0_12, output_MAC_0_13, output_MAC_0_14, output_MAC_0_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_1_0, output_MAC_1_1, output_MAC_1_2, output_MAC_1_3, output_MAC_1_4, output_MAC_1_5, output_MAC_1_6, output_MAC_1_7, output_MAC_1_8, output_MAC_1_9, 
		output_MAC_1_10, output_MAC_1_11, output_MAC_1_12, output_MAC_1_13, output_MAC_1_14, output_MAC_1_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_2_0, output_MAC_2_1, output_MAC_2_2, output_MAC_2_3, output_MAC_2_4, output_MAC_2_5, output_MAC_2_6, output_MAC_2_7, output_MAC_2_8, output_MAC_2_9, 
		output_MAC_2_10, output_MAC_2_11, output_MAC_2_12, output_MAC_2_13, output_MAC_2_14, output_MAC_2_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_3_0, output_MAC_3_1, output_MAC_3_2, output_MAC_3_3, output_MAC_3_4, output_MAC_3_5, output_MAC_3_6, output_MAC_3_7, output_MAC_3_8, output_MAC_3_9, 
		output_MAC_3_10, output_MAC_3_11, output_MAC_3_12, output_MAC_3_13, output_MAC_3_14, output_MAC_3_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_4_0, output_MAC_4_1, output_MAC_4_2, output_MAC_4_3, output_MAC_4_4, output_MAC_4_5, output_MAC_4_6, output_MAC_4_7, output_MAC_4_8, output_MAC_4_9, 
		output_MAC_4_10, output_MAC_4_11, output_MAC_4_12, output_MAC_4_13, output_MAC_4_14, output_MAC_4_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_5_0, output_MAC_5_1, output_MAC_5_2, output_MAC_5_3, output_MAC_5_4, output_MAC_5_5, output_MAC_5_6, output_MAC_5_7, output_MAC_5_8, output_MAC_5_9, 
		output_MAC_5_10, output_MAC_5_11, output_MAC_5_12, output_MAC_5_13, output_MAC_5_14, output_MAC_5_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_6_0, output_MAC_6_1, output_MAC_6_2, output_MAC_6_3, output_MAC_6_4, output_MAC_6_5, output_MAC_6_6, output_MAC_6_7, output_MAC_6_8, output_MAC_6_9, 
		output_MAC_6_10, output_MAC_6_11, output_MAC_6_12, output_MAC_6_13, output_MAC_6_14, output_MAC_6_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_7_0, output_MAC_7_1, output_MAC_7_2, output_MAC_7_3, output_MAC_7_4, output_MAC_7_5, output_MAC_7_6, output_MAC_7_7, output_MAC_7_8, output_MAC_7_9, 
		output_MAC_7_10, output_MAC_7_11, output_MAC_7_12, output_MAC_7_13, output_MAC_7_14, output_MAC_7_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_8_0, output_MAC_8_1, output_MAC_8_2, output_MAC_8_3, output_MAC_8_4, output_MAC_8_5, output_MAC_8_6, output_MAC_8_7, output_MAC_8_8, output_MAC_8_9, 
		output_MAC_8_10, output_MAC_8_11, output_MAC_8_12, output_MAC_8_13, output_MAC_8_14, output_MAC_8_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_9_0, output_MAC_9_1, output_MAC_9_2, output_MAC_9_3, output_MAC_9_4, output_MAC_9_5, output_MAC_9_6, output_MAC_9_7, output_MAC_9_8, output_MAC_9_9, 
		output_MAC_9_10, output_MAC_9_11, output_MAC_9_12, output_MAC_9_13, output_MAC_9_14, output_MAC_9_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_10_0, output_MAC_10_1, output_MAC_10_2, output_MAC_10_3, output_MAC_10_4, output_MAC_10_5, output_MAC_10_6, output_MAC_10_7, output_MAC_10_8, output_MAC_10_9, 
		output_MAC_10_10, output_MAC_10_11, output_MAC_10_12, output_MAC_10_13, output_MAC_10_14, output_MAC_10_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_11_0, output_MAC_11_1, output_MAC_11_2, output_MAC_11_3, output_MAC_11_4, output_MAC_11_5, output_MAC_11_6, output_MAC_11_7, output_MAC_11_8, output_MAC_11_9, 
		output_MAC_11_10, output_MAC_11_11, output_MAC_11_12, output_MAC_11_13, output_MAC_11_14, output_MAC_11_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_12_0, output_MAC_12_1, output_MAC_12_2, output_MAC_12_3, output_MAC_12_4, output_MAC_12_5, output_MAC_12_6, output_MAC_12_7, output_MAC_12_8, output_MAC_12_9, 
		output_MAC_12_10, output_MAC_12_11, output_MAC_12_12, output_MAC_12_13, output_MAC_12_14, output_MAC_12_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_13_0, output_MAC_13_1, output_MAC_13_2, output_MAC_13_3, output_MAC_13_4, output_MAC_13_5, output_MAC_13_6, output_MAC_13_7, output_MAC_13_8, output_MAC_13_9, 
		output_MAC_13_10, output_MAC_13_11, output_MAC_13_12, output_MAC_13_13, output_MAC_13_14, output_MAC_13_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_14_0, output_MAC_14_1, output_MAC_14_2, output_MAC_14_3, output_MAC_14_4, output_MAC_14_5, output_MAC_14_6, output_MAC_14_7, output_MAC_14_8, output_MAC_14_9, 
		output_MAC_14_10, output_MAC_14_11, output_MAC_14_12, output_MAC_14_13, output_MAC_14_14, output_MAC_14_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_15_0, output_MAC_15_1, output_MAC_15_2, output_MAC_15_3, output_MAC_15_4, output_MAC_15_5, output_MAC_15_6, output_MAC_15_7, output_MAC_15_8, output_MAC_15_9, 
		output_MAC_15_10, output_MAC_15_11, output_MAC_15_12, output_MAC_15_13, output_MAC_15_14, output_MAC_15_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_16_0, output_MAC_16_1, output_MAC_16_2, output_MAC_16_3, output_MAC_16_4, output_MAC_16_5, output_MAC_16_6, output_MAC_16_7, output_MAC_16_8, output_MAC_16_9, 
		output_MAC_16_10, output_MAC_16_11, output_MAC_16_12, output_MAC_16_13, output_MAC_16_14, output_MAC_16_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_17_0, output_MAC_17_1, output_MAC_17_2, output_MAC_17_3, output_MAC_17_4, output_MAC_17_5, output_MAC_17_6, output_MAC_17_7, output_MAC_17_8, output_MAC_17_9, 
		output_MAC_17_10, output_MAC_17_11, output_MAC_17_12, output_MAC_17_13, output_MAC_17_14, output_MAC_17_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_18_0, output_MAC_18_1, output_MAC_18_2, output_MAC_18_3, output_MAC_18_4, output_MAC_18_5, output_MAC_18_6, output_MAC_18_7, output_MAC_18_8, output_MAC_18_9, 
		output_MAC_18_10, output_MAC_18_11, output_MAC_18_12, output_MAC_18_13, output_MAC_18_14, output_MAC_18_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_19_0, output_MAC_19_1, output_MAC_19_2, output_MAC_19_3, output_MAC_19_4, output_MAC_19_5, output_MAC_19_6, output_MAC_19_7, output_MAC_19_8, output_MAC_19_9, 
		output_MAC_19_10, output_MAC_19_11, output_MAC_19_12, output_MAC_19_13, output_MAC_19_14, output_MAC_19_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_20_0, output_MAC_20_1, output_MAC_20_2, output_MAC_20_3, output_MAC_20_4, output_MAC_20_5, output_MAC_20_6, output_MAC_20_7, output_MAC_20_8, output_MAC_20_9, 
		output_MAC_20_10, output_MAC_20_11, output_MAC_20_12, output_MAC_20_13, output_MAC_20_14, output_MAC_20_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_21_0, output_MAC_21_1, output_MAC_21_2, output_MAC_21_3, output_MAC_21_4, output_MAC_21_5, output_MAC_21_6, output_MAC_21_7, output_MAC_21_8, output_MAC_21_9, 
		output_MAC_21_10, output_MAC_21_11, output_MAC_21_12, output_MAC_21_13, output_MAC_21_14, output_MAC_21_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_22_0, output_MAC_22_1, output_MAC_22_2, output_MAC_22_3, output_MAC_22_4, output_MAC_22_5, output_MAC_22_6, output_MAC_22_7, output_MAC_22_8, output_MAC_22_9, 
		output_MAC_22_10, output_MAC_22_11, output_MAC_22_12, output_MAC_22_13, output_MAC_22_14, output_MAC_22_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_23_0, output_MAC_23_1, output_MAC_23_2, output_MAC_23_3, output_MAC_23_4, output_MAC_23_5, output_MAC_23_6, output_MAC_23_7, output_MAC_23_8, output_MAC_23_9, 
		output_MAC_23_10, output_MAC_23_11, output_MAC_23_12, output_MAC_23_13, output_MAC_23_14, output_MAC_23_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_24_0, output_MAC_24_1, output_MAC_24_2, output_MAC_24_3, output_MAC_24_4, output_MAC_24_5, output_MAC_24_6, output_MAC_24_7, output_MAC_24_8, output_MAC_24_9, 
		output_MAC_24_10, output_MAC_24_11, output_MAC_24_12, output_MAC_24_13, output_MAC_24_14, output_MAC_24_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_25_0, output_MAC_25_1, output_MAC_25_2, output_MAC_25_3, output_MAC_25_4, output_MAC_25_5, output_MAC_25_6, output_MAC_25_7, output_MAC_25_8, output_MAC_25_9, 
		output_MAC_25_10, output_MAC_25_11, output_MAC_25_12, output_MAC_25_13, output_MAC_25_14, output_MAC_25_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_26_0, output_MAC_26_1, output_MAC_26_2, output_MAC_26_3, output_MAC_26_4, output_MAC_26_5, output_MAC_26_6, output_MAC_26_7, output_MAC_26_8, output_MAC_26_9, 
		output_MAC_26_10, output_MAC_26_11, output_MAC_26_12, output_MAC_26_13, output_MAC_26_14, output_MAC_26_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_27_0, output_MAC_27_1, output_MAC_27_2, output_MAC_27_3, output_MAC_27_4, output_MAC_27_5, output_MAC_27_6, output_MAC_27_7, output_MAC_27_8, output_MAC_27_9, 
		output_MAC_27_10, output_MAC_27_11, output_MAC_27_12, output_MAC_27_13, output_MAC_27_14, output_MAC_27_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_28_0, output_MAC_28_1, output_MAC_28_2, output_MAC_28_3, output_MAC_28_4, output_MAC_28_5, output_MAC_28_6, output_MAC_28_7, output_MAC_28_8, output_MAC_28_9, 
		output_MAC_28_10, output_MAC_28_11, output_MAC_28_12, output_MAC_28_13, output_MAC_28_14, output_MAC_28_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_29_0, output_MAC_29_1, output_MAC_29_2, output_MAC_29_3, output_MAC_29_4, output_MAC_29_5, output_MAC_29_6, output_MAC_29_7, output_MAC_29_8, output_MAC_29_9, 
		output_MAC_29_10, output_MAC_29_11, output_MAC_29_12, output_MAC_29_13, output_MAC_29_14, output_MAC_29_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_30_0, output_MAC_30_1, output_MAC_30_2, output_MAC_30_3, output_MAC_30_4, output_MAC_30_5, output_MAC_30_6, output_MAC_30_7, output_MAC_30_8, output_MAC_30_9, 
		output_MAC_30_10, output_MAC_30_11, output_MAC_30_12, output_MAC_30_13, output_MAC_30_14, output_MAC_30_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_31_0, output_MAC_31_1, output_MAC_31_2, output_MAC_31_3, output_MAC_31_4, output_MAC_31_5, output_MAC_31_6, output_MAC_31_7, output_MAC_31_8, output_MAC_31_9, 
		output_MAC_31_10, output_MAC_31_11, output_MAC_31_12, output_MAC_31_13, output_MAC_31_14, output_MAC_31_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_32_0, output_MAC_32_1, output_MAC_32_2, output_MAC_32_3, output_MAC_32_4, output_MAC_32_5, output_MAC_32_6, output_MAC_32_7, output_MAC_32_8, output_MAC_32_9, 
		output_MAC_32_10, output_MAC_32_11, output_MAC_32_12, output_MAC_32_13, output_MAC_32_14, output_MAC_32_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_33_0, output_MAC_33_1, output_MAC_33_2, output_MAC_33_3, output_MAC_33_4, output_MAC_33_5, output_MAC_33_6, output_MAC_33_7, output_MAC_33_8, output_MAC_33_9, 
		output_MAC_33_10, output_MAC_33_11, output_MAC_33_12, output_MAC_33_13, output_MAC_33_14, output_MAC_33_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_34_0, output_MAC_34_1, output_MAC_34_2, output_MAC_34_3, output_MAC_34_4, output_MAC_34_5, output_MAC_34_6, output_MAC_34_7, output_MAC_34_8, output_MAC_34_9, 
		output_MAC_34_10, output_MAC_34_11, output_MAC_34_12, output_MAC_34_13, output_MAC_34_14, output_MAC_34_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_35_0, output_MAC_35_1, output_MAC_35_2, output_MAC_35_3, output_MAC_35_4, output_MAC_35_5, output_MAC_35_6, output_MAC_35_7, output_MAC_35_8, output_MAC_35_9, 
		output_MAC_35_10, output_MAC_35_11, output_MAC_35_12, output_MAC_35_13, output_MAC_35_14, output_MAC_35_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_36_0, output_MAC_36_1, output_MAC_36_2, output_MAC_36_3, output_MAC_36_4, output_MAC_36_5, output_MAC_36_6, output_MAC_36_7, output_MAC_36_8, output_MAC_36_9, 
		output_MAC_36_10, output_MAC_36_11, output_MAC_36_12, output_MAC_36_13, output_MAC_36_14, output_MAC_36_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_37_0, output_MAC_37_1, output_MAC_37_2, output_MAC_37_3, output_MAC_37_4, output_MAC_37_5, output_MAC_37_6, output_MAC_37_7, output_MAC_37_8, output_MAC_37_9, 
		output_MAC_37_10, output_MAC_37_11, output_MAC_37_12, output_MAC_37_13, output_MAC_37_14, output_MAC_37_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_38_0, output_MAC_38_1, output_MAC_38_2, output_MAC_38_3, output_MAC_38_4, output_MAC_38_5, output_MAC_38_6, output_MAC_38_7, output_MAC_38_8, output_MAC_38_9, 
		output_MAC_38_10, output_MAC_38_11, output_MAC_38_12, output_MAC_38_13, output_MAC_38_14, output_MAC_38_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_39_0, output_MAC_39_1, output_MAC_39_2, output_MAC_39_3, output_MAC_39_4, output_MAC_39_5, output_MAC_39_6, output_MAC_39_7, output_MAC_39_8, output_MAC_39_9, 
		output_MAC_39_10, output_MAC_39_11, output_MAC_39_12, output_MAC_39_13, output_MAC_39_14, output_MAC_39_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_40_0, output_MAC_40_1, output_MAC_40_2, output_MAC_40_3, output_MAC_40_4, output_MAC_40_5, output_MAC_40_6, output_MAC_40_7, output_MAC_40_8, output_MAC_40_9, 
		output_MAC_40_10, output_MAC_40_11, output_MAC_40_12, output_MAC_40_13, output_MAC_40_14, output_MAC_40_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_41_0, output_MAC_41_1, output_MAC_41_2, output_MAC_41_3, output_MAC_41_4, output_MAC_41_5, output_MAC_41_6, output_MAC_41_7, output_MAC_41_8, output_MAC_41_9, 
		output_MAC_41_10, output_MAC_41_11, output_MAC_41_12, output_MAC_41_13, output_MAC_41_14, output_MAC_41_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_42_0, output_MAC_42_1, output_MAC_42_2, output_MAC_42_3, output_MAC_42_4, output_MAC_42_5, output_MAC_42_6, output_MAC_42_7, output_MAC_42_8, output_MAC_42_9, 
		output_MAC_42_10, output_MAC_42_11, output_MAC_42_12, output_MAC_42_13, output_MAC_42_14, output_MAC_42_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_43_0, output_MAC_43_1, output_MAC_43_2, output_MAC_43_3, output_MAC_43_4, output_MAC_43_5, output_MAC_43_6, output_MAC_43_7, output_MAC_43_8, output_MAC_43_9, 
		output_MAC_43_10, output_MAC_43_11, output_MAC_43_12, output_MAC_43_13, output_MAC_43_14, output_MAC_43_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_44_0, output_MAC_44_1, output_MAC_44_2, output_MAC_44_3, output_MAC_44_4, output_MAC_44_5, output_MAC_44_6, output_MAC_44_7, output_MAC_44_8, output_MAC_44_9, 
		output_MAC_44_10, output_MAC_44_11, output_MAC_44_12, output_MAC_44_13, output_MAC_44_14, output_MAC_44_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_45_0, output_MAC_45_1, output_MAC_45_2, output_MAC_45_3, output_MAC_45_4, output_MAC_45_5, output_MAC_45_6, output_MAC_45_7, output_MAC_45_8, output_MAC_45_9, 
		output_MAC_45_10, output_MAC_45_11, output_MAC_45_12, output_MAC_45_13, output_MAC_45_14, output_MAC_45_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_46_0, output_MAC_46_1, output_MAC_46_2, output_MAC_46_3, output_MAC_46_4, output_MAC_46_5, output_MAC_46_6, output_MAC_46_7, output_MAC_46_8, output_MAC_46_9, 
		output_MAC_46_10, output_MAC_46_11, output_MAC_46_12, output_MAC_46_13, output_MAC_46_14, output_MAC_46_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_47_0, output_MAC_47_1, output_MAC_47_2, output_MAC_47_3, output_MAC_47_4, output_MAC_47_5, output_MAC_47_6, output_MAC_47_7, output_MAC_47_8, output_MAC_47_9, 
		output_MAC_47_10, output_MAC_47_11, output_MAC_47_12, output_MAC_47_13, output_MAC_47_14, output_MAC_47_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_48_0, output_MAC_48_1, output_MAC_48_2, output_MAC_48_3, output_MAC_48_4, output_MAC_48_5, output_MAC_48_6, output_MAC_48_7, output_MAC_48_8, output_MAC_48_9, 
		output_MAC_48_10, output_MAC_48_11, output_MAC_48_12, output_MAC_48_13, output_MAC_48_14, output_MAC_48_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_49_0, output_MAC_49_1, output_MAC_49_2, output_MAC_49_3, output_MAC_49_4, output_MAC_49_5, output_MAC_49_6, output_MAC_49_7, output_MAC_49_8, output_MAC_49_9, 
		output_MAC_49_10, output_MAC_49_11, output_MAC_49_12, output_MAC_49_13, output_MAC_49_14, output_MAC_49_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_50_0, output_MAC_50_1, output_MAC_50_2, output_MAC_50_3, output_MAC_50_4, output_MAC_50_5, output_MAC_50_6, output_MAC_50_7, output_MAC_50_8, output_MAC_50_9, 
		output_MAC_50_10, output_MAC_50_11, output_MAC_50_12, output_MAC_50_13, output_MAC_50_14, output_MAC_50_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_51_0, output_MAC_51_1, output_MAC_51_2, output_MAC_51_3, output_MAC_51_4, output_MAC_51_5, output_MAC_51_6, output_MAC_51_7, output_MAC_51_8, output_MAC_51_9, 
		output_MAC_51_10, output_MAC_51_11, output_MAC_51_12, output_MAC_51_13, output_MAC_51_14, output_MAC_51_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_52_0, output_MAC_52_1, output_MAC_52_2, output_MAC_52_3, output_MAC_52_4, output_MAC_52_5, output_MAC_52_6, output_MAC_52_7, output_MAC_52_8, output_MAC_52_9, 
		output_MAC_52_10, output_MAC_52_11, output_MAC_52_12, output_MAC_52_13, output_MAC_52_14, output_MAC_52_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_53_0, output_MAC_53_1, output_MAC_53_2, output_MAC_53_3, output_MAC_53_4, output_MAC_53_5, output_MAC_53_6, output_MAC_53_7, output_MAC_53_8, output_MAC_53_9, 
		output_MAC_53_10, output_MAC_53_11, output_MAC_53_12, output_MAC_53_13, output_MAC_53_14, output_MAC_53_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_54_0, output_MAC_54_1, output_MAC_54_2, output_MAC_54_3, output_MAC_54_4, output_MAC_54_5, output_MAC_54_6, output_MAC_54_7, output_MAC_54_8, output_MAC_54_9, 
		output_MAC_54_10, output_MAC_54_11, output_MAC_54_12, output_MAC_54_13, output_MAC_54_14, output_MAC_54_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_55_0, output_MAC_55_1, output_MAC_55_2, output_MAC_55_3, output_MAC_55_4, output_MAC_55_5, output_MAC_55_6, output_MAC_55_7, output_MAC_55_8, output_MAC_55_9, 
		output_MAC_55_10, output_MAC_55_11, output_MAC_55_12, output_MAC_55_13, output_MAC_55_14, output_MAC_55_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_56_0, output_MAC_56_1, output_MAC_56_2, output_MAC_56_3, output_MAC_56_4, output_MAC_56_5, output_MAC_56_6, output_MAC_56_7, output_MAC_56_8, output_MAC_56_9, 
		output_MAC_56_10, output_MAC_56_11, output_MAC_56_12, output_MAC_56_13, output_MAC_56_14, output_MAC_56_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_57_0, output_MAC_57_1, output_MAC_57_2, output_MAC_57_3, output_MAC_57_4, output_MAC_57_5, output_MAC_57_6, output_MAC_57_7, output_MAC_57_8, output_MAC_57_9, 
		output_MAC_57_10, output_MAC_57_11, output_MAC_57_12, output_MAC_57_13, output_MAC_57_14, output_MAC_57_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_58_0, output_MAC_58_1, output_MAC_58_2, output_MAC_58_3, output_MAC_58_4, output_MAC_58_5, output_MAC_58_6, output_MAC_58_7, output_MAC_58_8, output_MAC_58_9, 
		output_MAC_58_10, output_MAC_58_11, output_MAC_58_12, output_MAC_58_13, output_MAC_58_14, output_MAC_58_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_59_0, output_MAC_59_1, output_MAC_59_2, output_MAC_59_3, output_MAC_59_4, output_MAC_59_5, output_MAC_59_6, output_MAC_59_7, output_MAC_59_8, output_MAC_59_9, 
		output_MAC_59_10, output_MAC_59_11, output_MAC_59_12, output_MAC_59_13, output_MAC_59_14, output_MAC_59_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_60_0, output_MAC_60_1, output_MAC_60_2, output_MAC_60_3, output_MAC_60_4, output_MAC_60_5, output_MAC_60_6, output_MAC_60_7, output_MAC_60_8, output_MAC_60_9, 
		output_MAC_60_10, output_MAC_60_11, output_MAC_60_12, output_MAC_60_13, output_MAC_60_14, output_MAC_60_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_61_0, output_MAC_61_1, output_MAC_61_2, output_MAC_61_3, output_MAC_61_4, output_MAC_61_5, output_MAC_61_6, output_MAC_61_7, output_MAC_61_8, output_MAC_61_9, 
		output_MAC_61_10, output_MAC_61_11, output_MAC_61_12, output_MAC_61_13, output_MAC_61_14, output_MAC_61_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_62_0, output_MAC_62_1, output_MAC_62_2, output_MAC_62_3, output_MAC_62_4, output_MAC_62_5, output_MAC_62_6, output_MAC_62_7, output_MAC_62_8, output_MAC_62_9, 
		output_MAC_62_10, output_MAC_62_11, output_MAC_62_12, output_MAC_62_13, output_MAC_62_14, output_MAC_62_15: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_63_0, output_MAC_63_1, output_MAC_63_2, output_MAC_63_3, output_MAC_63_4, output_MAC_63_5, output_MAC_63_6, output_MAC_63_7, output_MAC_63_8, output_MAC_63_9, 
		output_MAC_63_10, output_MAC_63_11, output_MAC_63_12, output_MAC_63_13, output_MAC_63_14, output_MAC_63_15: STD_LOGIC_VECTOR(31 downto 0);

BEGIN

	MAC_0_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_0, data_out=>output_MAC_0_0);
	MAC_0_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_1, data_out=>output_MAC_0_1);
	MAC_0_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_2, data_out=>output_MAC_0_2);
	MAC_0_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_3, data_out=>output_MAC_0_3);
	MAC_0_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_4, data_out=>output_MAC_0_4);
	MAC_0_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_5, data_out=>output_MAC_0_5);
	MAC_0_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_6, data_out=>output_MAC_0_6);
	MAC_0_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_7, data_out=>output_MAC_0_7);
	MAC_0_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_8, data_out=>output_MAC_0_8);
	MAC_0_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_9, data_out=>output_MAC_0_9);
	MAC_0_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_10, data_out=>output_MAC_0_10);
	MAC_0_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_11, data_out=>output_MAC_0_11);
	MAC_0_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_12, data_out=>output_MAC_0_12);
	MAC_0_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_13, data_out=>output_MAC_0_13);
	MAC_0_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_14, data_out=>output_MAC_0_14);
	MAC_0_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_15, data_out=>output_MAC_0_15);
	MAC_1_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_0, data_out=>output_MAC_1_0);
	MAC_1_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_1, data_out=>output_MAC_1_1);
	MAC_1_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_2, data_out=>output_MAC_1_2);
	MAC_1_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_3, data_out=>output_MAC_1_3);
	MAC_1_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_4, data_out=>output_MAC_1_4);
	MAC_1_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_5, data_out=>output_MAC_1_5);
	MAC_1_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_6, data_out=>output_MAC_1_6);
	MAC_1_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_7, data_out=>output_MAC_1_7);
	MAC_1_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_8, data_out=>output_MAC_1_8);
	MAC_1_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_9, data_out=>output_MAC_1_9);
	MAC_1_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_10, data_out=>output_MAC_1_10);
	MAC_1_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_11, data_out=>output_MAC_1_11);
	MAC_1_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_12, data_out=>output_MAC_1_12);
	MAC_1_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_13, data_out=>output_MAC_1_13);
	MAC_1_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_14, data_out=>output_MAC_1_14);
	MAC_1_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_15, data_out=>output_MAC_1_15);
	MAC_2_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_0, data_out=>output_MAC_2_0);
	MAC_2_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_1, data_out=>output_MAC_2_1);
	MAC_2_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_2, data_out=>output_MAC_2_2);
	MAC_2_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_3, data_out=>output_MAC_2_3);
	MAC_2_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_4, data_out=>output_MAC_2_4);
	MAC_2_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_5, data_out=>output_MAC_2_5);
	MAC_2_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_6, data_out=>output_MAC_2_6);
	MAC_2_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_7, data_out=>output_MAC_2_7);
	MAC_2_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_8, data_out=>output_MAC_2_8);
	MAC_2_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_9, data_out=>output_MAC_2_9);
	MAC_2_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_10, data_out=>output_MAC_2_10);
	MAC_2_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_11, data_out=>output_MAC_2_11);
	MAC_2_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_12, data_out=>output_MAC_2_12);
	MAC_2_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_13, data_out=>output_MAC_2_13);
	MAC_2_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_14, data_out=>output_MAC_2_14);
	MAC_2_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_15, data_out=>output_MAC_2_15);
	MAC_3_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_0, data_out=>output_MAC_3_0);
	MAC_3_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_1, data_out=>output_MAC_3_1);
	MAC_3_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_2, data_out=>output_MAC_3_2);
	MAC_3_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_3, data_out=>output_MAC_3_3);
	MAC_3_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_4, data_out=>output_MAC_3_4);
	MAC_3_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_5, data_out=>output_MAC_3_5);
	MAC_3_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_6, data_out=>output_MAC_3_6);
	MAC_3_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_7, data_out=>output_MAC_3_7);
	MAC_3_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_8, data_out=>output_MAC_3_8);
	MAC_3_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_9, data_out=>output_MAC_3_9);
	MAC_3_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_10, data_out=>output_MAC_3_10);
	MAC_3_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_11, data_out=>output_MAC_3_11);
	MAC_3_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_12, data_out=>output_MAC_3_12);
	MAC_3_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_13, data_out=>output_MAC_3_13);
	MAC_3_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_14, data_out=>output_MAC_3_14);
	MAC_3_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_15, data_out=>output_MAC_3_15);
	MAC_4_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_0, data_out=>output_MAC_4_0);
	MAC_4_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_1, data_out=>output_MAC_4_1);
	MAC_4_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_2, data_out=>output_MAC_4_2);
	MAC_4_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_3, data_out=>output_MAC_4_3);
	MAC_4_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_4, data_out=>output_MAC_4_4);
	MAC_4_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_5, data_out=>output_MAC_4_5);
	MAC_4_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_6, data_out=>output_MAC_4_6);
	MAC_4_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_7, data_out=>output_MAC_4_7);
	MAC_4_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_8, data_out=>output_MAC_4_8);
	MAC_4_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_9, data_out=>output_MAC_4_9);
	MAC_4_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_10, data_out=>output_MAC_4_10);
	MAC_4_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_11, data_out=>output_MAC_4_11);
	MAC_4_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_12, data_out=>output_MAC_4_12);
	MAC_4_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_13, data_out=>output_MAC_4_13);
	MAC_4_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_14, data_out=>output_MAC_4_14);
	MAC_4_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_15, data_out=>output_MAC_4_15);
	MAC_5_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_0, data_out=>output_MAC_5_0);
	MAC_5_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_1, data_out=>output_MAC_5_1);
	MAC_5_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_2, data_out=>output_MAC_5_2);
	MAC_5_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_3, data_out=>output_MAC_5_3);
	MAC_5_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_4, data_out=>output_MAC_5_4);
	MAC_5_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_5, data_out=>output_MAC_5_5);
	MAC_5_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_6, data_out=>output_MAC_5_6);
	MAC_5_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_7, data_out=>output_MAC_5_7);
	MAC_5_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_8, data_out=>output_MAC_5_8);
	MAC_5_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_9, data_out=>output_MAC_5_9);
	MAC_5_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_10, data_out=>output_MAC_5_10);
	MAC_5_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_11, data_out=>output_MAC_5_11);
	MAC_5_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_12, data_out=>output_MAC_5_12);
	MAC_5_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_13, data_out=>output_MAC_5_13);
	MAC_5_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_14, data_out=>output_MAC_5_14);
	MAC_5_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_15, data_out=>output_MAC_5_15);
	MAC_6_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_0, data_out=>output_MAC_6_0);
	MAC_6_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_1, data_out=>output_MAC_6_1);
	MAC_6_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_2, data_out=>output_MAC_6_2);
	MAC_6_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_3, data_out=>output_MAC_6_3);
	MAC_6_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_4, data_out=>output_MAC_6_4);
	MAC_6_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_5, data_out=>output_MAC_6_5);
	MAC_6_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_6, data_out=>output_MAC_6_6);
	MAC_6_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_7, data_out=>output_MAC_6_7);
	MAC_6_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_8, data_out=>output_MAC_6_8);
	MAC_6_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_9, data_out=>output_MAC_6_9);
	MAC_6_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_10, data_out=>output_MAC_6_10);
	MAC_6_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_11, data_out=>output_MAC_6_11);
	MAC_6_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_12, data_out=>output_MAC_6_12);
	MAC_6_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_13, data_out=>output_MAC_6_13);
	MAC_6_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_14, data_out=>output_MAC_6_14);
	MAC_6_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_15, data_out=>output_MAC_6_15);
	MAC_7_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_0, data_out=>output_MAC_7_0);
	MAC_7_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_1, data_out=>output_MAC_7_1);
	MAC_7_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_2, data_out=>output_MAC_7_2);
	MAC_7_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_3, data_out=>output_MAC_7_3);
	MAC_7_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_4, data_out=>output_MAC_7_4);
	MAC_7_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_5, data_out=>output_MAC_7_5);
	MAC_7_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_6, data_out=>output_MAC_7_6);
	MAC_7_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_7, data_out=>output_MAC_7_7);
	MAC_7_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_8, data_out=>output_MAC_7_8);
	MAC_7_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_9, data_out=>output_MAC_7_9);
	MAC_7_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_10, data_out=>output_MAC_7_10);
	MAC_7_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_11, data_out=>output_MAC_7_11);
	MAC_7_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_12, data_out=>output_MAC_7_12);
	MAC_7_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_13, data_out=>output_MAC_7_13);
	MAC_7_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_14, data_out=>output_MAC_7_14);
	MAC_7_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_15, data_out=>output_MAC_7_15);
	MAC_8_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_0, data_out=>output_MAC_8_0);
	MAC_8_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_1, data_out=>output_MAC_8_1);
	MAC_8_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_2, data_out=>output_MAC_8_2);
	MAC_8_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_3, data_out=>output_MAC_8_3);
	MAC_8_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_4, data_out=>output_MAC_8_4);
	MAC_8_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_5, data_out=>output_MAC_8_5);
	MAC_8_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_6, data_out=>output_MAC_8_6);
	MAC_8_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_7, data_out=>output_MAC_8_7);
	MAC_8_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_8, data_out=>output_MAC_8_8);
	MAC_8_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_9, data_out=>output_MAC_8_9);
	MAC_8_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_10, data_out=>output_MAC_8_10);
	MAC_8_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_11, data_out=>output_MAC_8_11);
	MAC_8_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_12, data_out=>output_MAC_8_12);
	MAC_8_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_13, data_out=>output_MAC_8_13);
	MAC_8_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_14, data_out=>output_MAC_8_14);
	MAC_8_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_8, data_in_B=>input_col_15, data_out=>output_MAC_8_15);
	MAC_9_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_0, data_out=>output_MAC_9_0);
	MAC_9_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_1, data_out=>output_MAC_9_1);
	MAC_9_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_2, data_out=>output_MAC_9_2);
	MAC_9_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_3, data_out=>output_MAC_9_3);
	MAC_9_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_4, data_out=>output_MAC_9_4);
	MAC_9_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_5, data_out=>output_MAC_9_5);
	MAC_9_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_6, data_out=>output_MAC_9_6);
	MAC_9_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_7, data_out=>output_MAC_9_7);
	MAC_9_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_8, data_out=>output_MAC_9_8);
	MAC_9_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_9, data_out=>output_MAC_9_9);
	MAC_9_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_10, data_out=>output_MAC_9_10);
	MAC_9_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_11, data_out=>output_MAC_9_11);
	MAC_9_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_12, data_out=>output_MAC_9_12);
	MAC_9_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_13, data_out=>output_MAC_9_13);
	MAC_9_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_14, data_out=>output_MAC_9_14);
	MAC_9_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_9, data_in_B=>input_col_15, data_out=>output_MAC_9_15);
	MAC_10_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_0, data_out=>output_MAC_10_0);
	MAC_10_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_1, data_out=>output_MAC_10_1);
	MAC_10_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_2, data_out=>output_MAC_10_2);
	MAC_10_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_3, data_out=>output_MAC_10_3);
	MAC_10_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_4, data_out=>output_MAC_10_4);
	MAC_10_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_5, data_out=>output_MAC_10_5);
	MAC_10_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_6, data_out=>output_MAC_10_6);
	MAC_10_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_7, data_out=>output_MAC_10_7);
	MAC_10_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_8, data_out=>output_MAC_10_8);
	MAC_10_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_9, data_out=>output_MAC_10_9);
	MAC_10_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_10, data_out=>output_MAC_10_10);
	MAC_10_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_11, data_out=>output_MAC_10_11);
	MAC_10_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_12, data_out=>output_MAC_10_12);
	MAC_10_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_13, data_out=>output_MAC_10_13);
	MAC_10_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_14, data_out=>output_MAC_10_14);
	MAC_10_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_10, data_in_B=>input_col_15, data_out=>output_MAC_10_15);
	MAC_11_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_0, data_out=>output_MAC_11_0);
	MAC_11_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_1, data_out=>output_MAC_11_1);
	MAC_11_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_2, data_out=>output_MAC_11_2);
	MAC_11_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_3, data_out=>output_MAC_11_3);
	MAC_11_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_4, data_out=>output_MAC_11_4);
	MAC_11_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_5, data_out=>output_MAC_11_5);
	MAC_11_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_6, data_out=>output_MAC_11_6);
	MAC_11_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_7, data_out=>output_MAC_11_7);
	MAC_11_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_8, data_out=>output_MAC_11_8);
	MAC_11_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_9, data_out=>output_MAC_11_9);
	MAC_11_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_10, data_out=>output_MAC_11_10);
	MAC_11_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_11, data_out=>output_MAC_11_11);
	MAC_11_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_12, data_out=>output_MAC_11_12);
	MAC_11_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_13, data_out=>output_MAC_11_13);
	MAC_11_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_14, data_out=>output_MAC_11_14);
	MAC_11_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_11, data_in_B=>input_col_15, data_out=>output_MAC_11_15);
	MAC_12_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_0, data_out=>output_MAC_12_0);
	MAC_12_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_1, data_out=>output_MAC_12_1);
	MAC_12_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_2, data_out=>output_MAC_12_2);
	MAC_12_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_3, data_out=>output_MAC_12_3);
	MAC_12_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_4, data_out=>output_MAC_12_4);
	MAC_12_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_5, data_out=>output_MAC_12_5);
	MAC_12_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_6, data_out=>output_MAC_12_6);
	MAC_12_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_7, data_out=>output_MAC_12_7);
	MAC_12_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_8, data_out=>output_MAC_12_8);
	MAC_12_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_9, data_out=>output_MAC_12_9);
	MAC_12_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_10, data_out=>output_MAC_12_10);
	MAC_12_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_11, data_out=>output_MAC_12_11);
	MAC_12_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_12, data_out=>output_MAC_12_12);
	MAC_12_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_13, data_out=>output_MAC_12_13);
	MAC_12_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_14, data_out=>output_MAC_12_14);
	MAC_12_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_12, data_in_B=>input_col_15, data_out=>output_MAC_12_15);
	MAC_13_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_0, data_out=>output_MAC_13_0);
	MAC_13_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_1, data_out=>output_MAC_13_1);
	MAC_13_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_2, data_out=>output_MAC_13_2);
	MAC_13_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_3, data_out=>output_MAC_13_3);
	MAC_13_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_4, data_out=>output_MAC_13_4);
	MAC_13_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_5, data_out=>output_MAC_13_5);
	MAC_13_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_6, data_out=>output_MAC_13_6);
	MAC_13_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_7, data_out=>output_MAC_13_7);
	MAC_13_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_8, data_out=>output_MAC_13_8);
	MAC_13_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_9, data_out=>output_MAC_13_9);
	MAC_13_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_10, data_out=>output_MAC_13_10);
	MAC_13_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_11, data_out=>output_MAC_13_11);
	MAC_13_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_12, data_out=>output_MAC_13_12);
	MAC_13_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_13, data_out=>output_MAC_13_13);
	MAC_13_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_14, data_out=>output_MAC_13_14);
	MAC_13_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_13, data_in_B=>input_col_15, data_out=>output_MAC_13_15);
	MAC_14_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_0, data_out=>output_MAC_14_0);
	MAC_14_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_1, data_out=>output_MAC_14_1);
	MAC_14_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_2, data_out=>output_MAC_14_2);
	MAC_14_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_3, data_out=>output_MAC_14_3);
	MAC_14_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_4, data_out=>output_MAC_14_4);
	MAC_14_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_5, data_out=>output_MAC_14_5);
	MAC_14_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_6, data_out=>output_MAC_14_6);
	MAC_14_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_7, data_out=>output_MAC_14_7);
	MAC_14_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_8, data_out=>output_MAC_14_8);
	MAC_14_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_9, data_out=>output_MAC_14_9);
	MAC_14_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_10, data_out=>output_MAC_14_10);
	MAC_14_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_11, data_out=>output_MAC_14_11);
	MAC_14_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_12, data_out=>output_MAC_14_12);
	MAC_14_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_13, data_out=>output_MAC_14_13);
	MAC_14_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_14, data_out=>output_MAC_14_14);
	MAC_14_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_14, data_in_B=>input_col_15, data_out=>output_MAC_14_15);
	MAC_15_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_0, data_out=>output_MAC_15_0);
	MAC_15_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_1, data_out=>output_MAC_15_1);
	MAC_15_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_2, data_out=>output_MAC_15_2);
	MAC_15_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_3, data_out=>output_MAC_15_3);
	MAC_15_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_4, data_out=>output_MAC_15_4);
	MAC_15_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_5, data_out=>output_MAC_15_5);
	MAC_15_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_6, data_out=>output_MAC_15_6);
	MAC_15_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_7, data_out=>output_MAC_15_7);
	MAC_15_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_8, data_out=>output_MAC_15_8);
	MAC_15_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_9, data_out=>output_MAC_15_9);
	MAC_15_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_10, data_out=>output_MAC_15_10);
	MAC_15_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_11, data_out=>output_MAC_15_11);
	MAC_15_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_12, data_out=>output_MAC_15_12);
	MAC_15_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_13, data_out=>output_MAC_15_13);
	MAC_15_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_14, data_out=>output_MAC_15_14);
	MAC_15_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_15, data_in_B=>input_col_15, data_out=>output_MAC_15_15);
	MAC_16_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_0, data_out=>output_MAC_16_0);
	MAC_16_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_1, data_out=>output_MAC_16_1);
	MAC_16_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_2, data_out=>output_MAC_16_2);
	MAC_16_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_3, data_out=>output_MAC_16_3);
	MAC_16_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_4, data_out=>output_MAC_16_4);
	MAC_16_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_5, data_out=>output_MAC_16_5);
	MAC_16_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_6, data_out=>output_MAC_16_6);
	MAC_16_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_7, data_out=>output_MAC_16_7);
	MAC_16_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_8, data_out=>output_MAC_16_8);
	MAC_16_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_9, data_out=>output_MAC_16_9);
	MAC_16_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_10, data_out=>output_MAC_16_10);
	MAC_16_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_11, data_out=>output_MAC_16_11);
	MAC_16_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_12, data_out=>output_MAC_16_12);
	MAC_16_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_13, data_out=>output_MAC_16_13);
	MAC_16_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_14, data_out=>output_MAC_16_14);
	MAC_16_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_16, data_in_B=>input_col_15, data_out=>output_MAC_16_15);
	MAC_17_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_0, data_out=>output_MAC_17_0);
	MAC_17_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_1, data_out=>output_MAC_17_1);
	MAC_17_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_2, data_out=>output_MAC_17_2);
	MAC_17_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_3, data_out=>output_MAC_17_3);
	MAC_17_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_4, data_out=>output_MAC_17_4);
	MAC_17_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_5, data_out=>output_MAC_17_5);
	MAC_17_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_6, data_out=>output_MAC_17_6);
	MAC_17_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_7, data_out=>output_MAC_17_7);
	MAC_17_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_8, data_out=>output_MAC_17_8);
	MAC_17_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_9, data_out=>output_MAC_17_9);
	MAC_17_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_10, data_out=>output_MAC_17_10);
	MAC_17_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_11, data_out=>output_MAC_17_11);
	MAC_17_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_12, data_out=>output_MAC_17_12);
	MAC_17_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_13, data_out=>output_MAC_17_13);
	MAC_17_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_14, data_out=>output_MAC_17_14);
	MAC_17_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_17, data_in_B=>input_col_15, data_out=>output_MAC_17_15);
	MAC_18_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_0, data_out=>output_MAC_18_0);
	MAC_18_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_1, data_out=>output_MAC_18_1);
	MAC_18_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_2, data_out=>output_MAC_18_2);
	MAC_18_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_3, data_out=>output_MAC_18_3);
	MAC_18_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_4, data_out=>output_MAC_18_4);
	MAC_18_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_5, data_out=>output_MAC_18_5);
	MAC_18_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_6, data_out=>output_MAC_18_6);
	MAC_18_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_7, data_out=>output_MAC_18_7);
	MAC_18_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_8, data_out=>output_MAC_18_8);
	MAC_18_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_9, data_out=>output_MAC_18_9);
	MAC_18_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_10, data_out=>output_MAC_18_10);
	MAC_18_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_11, data_out=>output_MAC_18_11);
	MAC_18_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_12, data_out=>output_MAC_18_12);
	MAC_18_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_13, data_out=>output_MAC_18_13);
	MAC_18_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_14, data_out=>output_MAC_18_14);
	MAC_18_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_18, data_in_B=>input_col_15, data_out=>output_MAC_18_15);
	MAC_19_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_0, data_out=>output_MAC_19_0);
	MAC_19_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_1, data_out=>output_MAC_19_1);
	MAC_19_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_2, data_out=>output_MAC_19_2);
	MAC_19_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_3, data_out=>output_MAC_19_3);
	MAC_19_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_4, data_out=>output_MAC_19_4);
	MAC_19_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_5, data_out=>output_MAC_19_5);
	MAC_19_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_6, data_out=>output_MAC_19_6);
	MAC_19_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_7, data_out=>output_MAC_19_7);
	MAC_19_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_8, data_out=>output_MAC_19_8);
	MAC_19_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_9, data_out=>output_MAC_19_9);
	MAC_19_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_10, data_out=>output_MAC_19_10);
	MAC_19_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_11, data_out=>output_MAC_19_11);
	MAC_19_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_12, data_out=>output_MAC_19_12);
	MAC_19_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_13, data_out=>output_MAC_19_13);
	MAC_19_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_14, data_out=>output_MAC_19_14);
	MAC_19_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_19, data_in_B=>input_col_15, data_out=>output_MAC_19_15);
	MAC_20_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_0, data_out=>output_MAC_20_0);
	MAC_20_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_1, data_out=>output_MAC_20_1);
	MAC_20_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_2, data_out=>output_MAC_20_2);
	MAC_20_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_3, data_out=>output_MAC_20_3);
	MAC_20_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_4, data_out=>output_MAC_20_4);
	MAC_20_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_5, data_out=>output_MAC_20_5);
	MAC_20_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_6, data_out=>output_MAC_20_6);
	MAC_20_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_7, data_out=>output_MAC_20_7);
	MAC_20_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_8, data_out=>output_MAC_20_8);
	MAC_20_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_9, data_out=>output_MAC_20_9);
	MAC_20_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_10, data_out=>output_MAC_20_10);
	MAC_20_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_11, data_out=>output_MAC_20_11);
	MAC_20_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_12, data_out=>output_MAC_20_12);
	MAC_20_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_13, data_out=>output_MAC_20_13);
	MAC_20_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_14, data_out=>output_MAC_20_14);
	MAC_20_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_20, data_in_B=>input_col_15, data_out=>output_MAC_20_15);
	MAC_21_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_0, data_out=>output_MAC_21_0);
	MAC_21_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_1, data_out=>output_MAC_21_1);
	MAC_21_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_2, data_out=>output_MAC_21_2);
	MAC_21_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_3, data_out=>output_MAC_21_3);
	MAC_21_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_4, data_out=>output_MAC_21_4);
	MAC_21_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_5, data_out=>output_MAC_21_5);
	MAC_21_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_6, data_out=>output_MAC_21_6);
	MAC_21_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_7, data_out=>output_MAC_21_7);
	MAC_21_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_8, data_out=>output_MAC_21_8);
	MAC_21_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_9, data_out=>output_MAC_21_9);
	MAC_21_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_10, data_out=>output_MAC_21_10);
	MAC_21_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_11, data_out=>output_MAC_21_11);
	MAC_21_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_12, data_out=>output_MAC_21_12);
	MAC_21_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_13, data_out=>output_MAC_21_13);
	MAC_21_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_14, data_out=>output_MAC_21_14);
	MAC_21_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_21, data_in_B=>input_col_15, data_out=>output_MAC_21_15);
	MAC_22_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_0, data_out=>output_MAC_22_0);
	MAC_22_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_1, data_out=>output_MAC_22_1);
	MAC_22_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_2, data_out=>output_MAC_22_2);
	MAC_22_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_3, data_out=>output_MAC_22_3);
	MAC_22_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_4, data_out=>output_MAC_22_4);
	MAC_22_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_5, data_out=>output_MAC_22_5);
	MAC_22_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_6, data_out=>output_MAC_22_6);
	MAC_22_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_7, data_out=>output_MAC_22_7);
	MAC_22_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_8, data_out=>output_MAC_22_8);
	MAC_22_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_9, data_out=>output_MAC_22_9);
	MAC_22_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_10, data_out=>output_MAC_22_10);
	MAC_22_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_11, data_out=>output_MAC_22_11);
	MAC_22_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_12, data_out=>output_MAC_22_12);
	MAC_22_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_13, data_out=>output_MAC_22_13);
	MAC_22_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_14, data_out=>output_MAC_22_14);
	MAC_22_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_22, data_in_B=>input_col_15, data_out=>output_MAC_22_15);
	MAC_23_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_0, data_out=>output_MAC_23_0);
	MAC_23_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_1, data_out=>output_MAC_23_1);
	MAC_23_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_2, data_out=>output_MAC_23_2);
	MAC_23_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_3, data_out=>output_MAC_23_3);
	MAC_23_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_4, data_out=>output_MAC_23_4);
	MAC_23_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_5, data_out=>output_MAC_23_5);
	MAC_23_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_6, data_out=>output_MAC_23_6);
	MAC_23_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_7, data_out=>output_MAC_23_7);
	MAC_23_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_8, data_out=>output_MAC_23_8);
	MAC_23_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_9, data_out=>output_MAC_23_9);
	MAC_23_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_10, data_out=>output_MAC_23_10);
	MAC_23_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_11, data_out=>output_MAC_23_11);
	MAC_23_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_12, data_out=>output_MAC_23_12);
	MAC_23_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_13, data_out=>output_MAC_23_13);
	MAC_23_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_14, data_out=>output_MAC_23_14);
	MAC_23_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_23, data_in_B=>input_col_15, data_out=>output_MAC_23_15);
	MAC_24_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_0, data_out=>output_MAC_24_0);
	MAC_24_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_1, data_out=>output_MAC_24_1);
	MAC_24_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_2, data_out=>output_MAC_24_2);
	MAC_24_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_3, data_out=>output_MAC_24_3);
	MAC_24_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_4, data_out=>output_MAC_24_4);
	MAC_24_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_5, data_out=>output_MAC_24_5);
	MAC_24_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_6, data_out=>output_MAC_24_6);
	MAC_24_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_7, data_out=>output_MAC_24_7);
	MAC_24_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_8, data_out=>output_MAC_24_8);
	MAC_24_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_9, data_out=>output_MAC_24_9);
	MAC_24_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_10, data_out=>output_MAC_24_10);
	MAC_24_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_11, data_out=>output_MAC_24_11);
	MAC_24_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_12, data_out=>output_MAC_24_12);
	MAC_24_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_13, data_out=>output_MAC_24_13);
	MAC_24_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_14, data_out=>output_MAC_24_14);
	MAC_24_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_24, data_in_B=>input_col_15, data_out=>output_MAC_24_15);
	MAC_25_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_0, data_out=>output_MAC_25_0);
	MAC_25_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_1, data_out=>output_MAC_25_1);
	MAC_25_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_2, data_out=>output_MAC_25_2);
	MAC_25_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_3, data_out=>output_MAC_25_3);
	MAC_25_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_4, data_out=>output_MAC_25_4);
	MAC_25_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_5, data_out=>output_MAC_25_5);
	MAC_25_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_6, data_out=>output_MAC_25_6);
	MAC_25_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_7, data_out=>output_MAC_25_7);
	MAC_25_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_8, data_out=>output_MAC_25_8);
	MAC_25_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_9, data_out=>output_MAC_25_9);
	MAC_25_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_10, data_out=>output_MAC_25_10);
	MAC_25_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_11, data_out=>output_MAC_25_11);
	MAC_25_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_12, data_out=>output_MAC_25_12);
	MAC_25_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_13, data_out=>output_MAC_25_13);
	MAC_25_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_14, data_out=>output_MAC_25_14);
	MAC_25_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_25, data_in_B=>input_col_15, data_out=>output_MAC_25_15);
	MAC_26_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_0, data_out=>output_MAC_26_0);
	MAC_26_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_1, data_out=>output_MAC_26_1);
	MAC_26_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_2, data_out=>output_MAC_26_2);
	MAC_26_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_3, data_out=>output_MAC_26_3);
	MAC_26_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_4, data_out=>output_MAC_26_4);
	MAC_26_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_5, data_out=>output_MAC_26_5);
	MAC_26_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_6, data_out=>output_MAC_26_6);
	MAC_26_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_7, data_out=>output_MAC_26_7);
	MAC_26_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_8, data_out=>output_MAC_26_8);
	MAC_26_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_9, data_out=>output_MAC_26_9);
	MAC_26_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_10, data_out=>output_MAC_26_10);
	MAC_26_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_11, data_out=>output_MAC_26_11);
	MAC_26_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_12, data_out=>output_MAC_26_12);
	MAC_26_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_13, data_out=>output_MAC_26_13);
	MAC_26_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_14, data_out=>output_MAC_26_14);
	MAC_26_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_26, data_in_B=>input_col_15, data_out=>output_MAC_26_15);
	MAC_27_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_0, data_out=>output_MAC_27_0);
	MAC_27_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_1, data_out=>output_MAC_27_1);
	MAC_27_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_2, data_out=>output_MAC_27_2);
	MAC_27_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_3, data_out=>output_MAC_27_3);
	MAC_27_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_4, data_out=>output_MAC_27_4);
	MAC_27_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_5, data_out=>output_MAC_27_5);
	MAC_27_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_6, data_out=>output_MAC_27_6);
	MAC_27_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_7, data_out=>output_MAC_27_7);
	MAC_27_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_8, data_out=>output_MAC_27_8);
	MAC_27_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_9, data_out=>output_MAC_27_9);
	MAC_27_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_10, data_out=>output_MAC_27_10);
	MAC_27_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_11, data_out=>output_MAC_27_11);
	MAC_27_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_12, data_out=>output_MAC_27_12);
	MAC_27_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_13, data_out=>output_MAC_27_13);
	MAC_27_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_14, data_out=>output_MAC_27_14);
	MAC_27_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_27, data_in_B=>input_col_15, data_out=>output_MAC_27_15);
	MAC_28_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_0, data_out=>output_MAC_28_0);
	MAC_28_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_1, data_out=>output_MAC_28_1);
	MAC_28_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_2, data_out=>output_MAC_28_2);
	MAC_28_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_3, data_out=>output_MAC_28_3);
	MAC_28_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_4, data_out=>output_MAC_28_4);
	MAC_28_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_5, data_out=>output_MAC_28_5);
	MAC_28_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_6, data_out=>output_MAC_28_6);
	MAC_28_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_7, data_out=>output_MAC_28_7);
	MAC_28_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_8, data_out=>output_MAC_28_8);
	MAC_28_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_9, data_out=>output_MAC_28_9);
	MAC_28_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_10, data_out=>output_MAC_28_10);
	MAC_28_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_11, data_out=>output_MAC_28_11);
	MAC_28_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_12, data_out=>output_MAC_28_12);
	MAC_28_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_13, data_out=>output_MAC_28_13);
	MAC_28_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_14, data_out=>output_MAC_28_14);
	MAC_28_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_28, data_in_B=>input_col_15, data_out=>output_MAC_28_15);
	MAC_29_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_0, data_out=>output_MAC_29_0);
	MAC_29_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_1, data_out=>output_MAC_29_1);
	MAC_29_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_2, data_out=>output_MAC_29_2);
	MAC_29_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_3, data_out=>output_MAC_29_3);
	MAC_29_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_4, data_out=>output_MAC_29_4);
	MAC_29_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_5, data_out=>output_MAC_29_5);
	MAC_29_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_6, data_out=>output_MAC_29_6);
	MAC_29_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_7, data_out=>output_MAC_29_7);
	MAC_29_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_8, data_out=>output_MAC_29_8);
	MAC_29_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_9, data_out=>output_MAC_29_9);
	MAC_29_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_10, data_out=>output_MAC_29_10);
	MAC_29_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_11, data_out=>output_MAC_29_11);
	MAC_29_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_12, data_out=>output_MAC_29_12);
	MAC_29_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_13, data_out=>output_MAC_29_13);
	MAC_29_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_14, data_out=>output_MAC_29_14);
	MAC_29_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_29, data_in_B=>input_col_15, data_out=>output_MAC_29_15);
	MAC_30_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_0, data_out=>output_MAC_30_0);
	MAC_30_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_1, data_out=>output_MAC_30_1);
	MAC_30_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_2, data_out=>output_MAC_30_2);
	MAC_30_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_3, data_out=>output_MAC_30_3);
	MAC_30_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_4, data_out=>output_MAC_30_4);
	MAC_30_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_5, data_out=>output_MAC_30_5);
	MAC_30_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_6, data_out=>output_MAC_30_6);
	MAC_30_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_7, data_out=>output_MAC_30_7);
	MAC_30_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_8, data_out=>output_MAC_30_8);
	MAC_30_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_9, data_out=>output_MAC_30_9);
	MAC_30_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_10, data_out=>output_MAC_30_10);
	MAC_30_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_11, data_out=>output_MAC_30_11);
	MAC_30_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_12, data_out=>output_MAC_30_12);
	MAC_30_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_13, data_out=>output_MAC_30_13);
	MAC_30_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_14, data_out=>output_MAC_30_14);
	MAC_30_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_30, data_in_B=>input_col_15, data_out=>output_MAC_30_15);
	MAC_31_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_0, data_out=>output_MAC_31_0);
	MAC_31_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_1, data_out=>output_MAC_31_1);
	MAC_31_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_2, data_out=>output_MAC_31_2);
	MAC_31_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_3, data_out=>output_MAC_31_3);
	MAC_31_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_4, data_out=>output_MAC_31_4);
	MAC_31_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_5, data_out=>output_MAC_31_5);
	MAC_31_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_6, data_out=>output_MAC_31_6);
	MAC_31_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_7, data_out=>output_MAC_31_7);
	MAC_31_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_8, data_out=>output_MAC_31_8);
	MAC_31_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_9, data_out=>output_MAC_31_9);
	MAC_31_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_10, data_out=>output_MAC_31_10);
	MAC_31_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_11, data_out=>output_MAC_31_11);
	MAC_31_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_12, data_out=>output_MAC_31_12);
	MAC_31_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_13, data_out=>output_MAC_31_13);
	MAC_31_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_14, data_out=>output_MAC_31_14);
	MAC_31_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_31, data_in_B=>input_col_15, data_out=>output_MAC_31_15);
	MAC_32_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_0, data_out=>output_MAC_32_0);
	MAC_32_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_1, data_out=>output_MAC_32_1);
	MAC_32_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_2, data_out=>output_MAC_32_2);
	MAC_32_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_3, data_out=>output_MAC_32_3);
	MAC_32_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_4, data_out=>output_MAC_32_4);
	MAC_32_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_5, data_out=>output_MAC_32_5);
	MAC_32_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_6, data_out=>output_MAC_32_6);
	MAC_32_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_7, data_out=>output_MAC_32_7);
	MAC_32_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_8, data_out=>output_MAC_32_8);
	MAC_32_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_9, data_out=>output_MAC_32_9);
	MAC_32_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_10, data_out=>output_MAC_32_10);
	MAC_32_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_11, data_out=>output_MAC_32_11);
	MAC_32_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_12, data_out=>output_MAC_32_12);
	MAC_32_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_13, data_out=>output_MAC_32_13);
	MAC_32_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_14, data_out=>output_MAC_32_14);
	MAC_32_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_32, data_in_B=>input_col_15, data_out=>output_MAC_32_15);
	MAC_33_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_0, data_out=>output_MAC_33_0);
	MAC_33_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_1, data_out=>output_MAC_33_1);
	MAC_33_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_2, data_out=>output_MAC_33_2);
	MAC_33_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_3, data_out=>output_MAC_33_3);
	MAC_33_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_4, data_out=>output_MAC_33_4);
	MAC_33_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_5, data_out=>output_MAC_33_5);
	MAC_33_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_6, data_out=>output_MAC_33_6);
	MAC_33_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_7, data_out=>output_MAC_33_7);
	MAC_33_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_8, data_out=>output_MAC_33_8);
	MAC_33_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_9, data_out=>output_MAC_33_9);
	MAC_33_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_10, data_out=>output_MAC_33_10);
	MAC_33_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_11, data_out=>output_MAC_33_11);
	MAC_33_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_12, data_out=>output_MAC_33_12);
	MAC_33_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_13, data_out=>output_MAC_33_13);
	MAC_33_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_14, data_out=>output_MAC_33_14);
	MAC_33_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_33, data_in_B=>input_col_15, data_out=>output_MAC_33_15);
	MAC_34_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_0, data_out=>output_MAC_34_0);
	MAC_34_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_1, data_out=>output_MAC_34_1);
	MAC_34_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_2, data_out=>output_MAC_34_2);
	MAC_34_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_3, data_out=>output_MAC_34_3);
	MAC_34_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_4, data_out=>output_MAC_34_4);
	MAC_34_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_5, data_out=>output_MAC_34_5);
	MAC_34_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_6, data_out=>output_MAC_34_6);
	MAC_34_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_7, data_out=>output_MAC_34_7);
	MAC_34_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_8, data_out=>output_MAC_34_8);
	MAC_34_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_9, data_out=>output_MAC_34_9);
	MAC_34_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_10, data_out=>output_MAC_34_10);
	MAC_34_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_11, data_out=>output_MAC_34_11);
	MAC_34_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_12, data_out=>output_MAC_34_12);
	MAC_34_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_13, data_out=>output_MAC_34_13);
	MAC_34_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_14, data_out=>output_MAC_34_14);
	MAC_34_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_34, data_in_B=>input_col_15, data_out=>output_MAC_34_15);
	MAC_35_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_0, data_out=>output_MAC_35_0);
	MAC_35_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_1, data_out=>output_MAC_35_1);
	MAC_35_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_2, data_out=>output_MAC_35_2);
	MAC_35_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_3, data_out=>output_MAC_35_3);
	MAC_35_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_4, data_out=>output_MAC_35_4);
	MAC_35_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_5, data_out=>output_MAC_35_5);
	MAC_35_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_6, data_out=>output_MAC_35_6);
	MAC_35_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_7, data_out=>output_MAC_35_7);
	MAC_35_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_8, data_out=>output_MAC_35_8);
	MAC_35_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_9, data_out=>output_MAC_35_9);
	MAC_35_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_10, data_out=>output_MAC_35_10);
	MAC_35_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_11, data_out=>output_MAC_35_11);
	MAC_35_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_12, data_out=>output_MAC_35_12);
	MAC_35_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_13, data_out=>output_MAC_35_13);
	MAC_35_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_14, data_out=>output_MAC_35_14);
	MAC_35_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_35, data_in_B=>input_col_15, data_out=>output_MAC_35_15);
	MAC_36_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_0, data_out=>output_MAC_36_0);
	MAC_36_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_1, data_out=>output_MAC_36_1);
	MAC_36_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_2, data_out=>output_MAC_36_2);
	MAC_36_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_3, data_out=>output_MAC_36_3);
	MAC_36_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_4, data_out=>output_MAC_36_4);
	MAC_36_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_5, data_out=>output_MAC_36_5);
	MAC_36_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_6, data_out=>output_MAC_36_6);
	MAC_36_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_7, data_out=>output_MAC_36_7);
	MAC_36_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_8, data_out=>output_MAC_36_8);
	MAC_36_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_9, data_out=>output_MAC_36_9);
	MAC_36_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_10, data_out=>output_MAC_36_10);
	MAC_36_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_11, data_out=>output_MAC_36_11);
	MAC_36_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_12, data_out=>output_MAC_36_12);
	MAC_36_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_13, data_out=>output_MAC_36_13);
	MAC_36_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_14, data_out=>output_MAC_36_14);
	MAC_36_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_36, data_in_B=>input_col_15, data_out=>output_MAC_36_15);
	MAC_37_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_0, data_out=>output_MAC_37_0);
	MAC_37_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_1, data_out=>output_MAC_37_1);
	MAC_37_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_2, data_out=>output_MAC_37_2);
	MAC_37_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_3, data_out=>output_MAC_37_3);
	MAC_37_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_4, data_out=>output_MAC_37_4);
	MAC_37_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_5, data_out=>output_MAC_37_5);
	MAC_37_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_6, data_out=>output_MAC_37_6);
	MAC_37_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_7, data_out=>output_MAC_37_7);
	MAC_37_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_8, data_out=>output_MAC_37_8);
	MAC_37_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_9, data_out=>output_MAC_37_9);
	MAC_37_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_10, data_out=>output_MAC_37_10);
	MAC_37_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_11, data_out=>output_MAC_37_11);
	MAC_37_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_12, data_out=>output_MAC_37_12);
	MAC_37_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_13, data_out=>output_MAC_37_13);
	MAC_37_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_14, data_out=>output_MAC_37_14);
	MAC_37_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_37, data_in_B=>input_col_15, data_out=>output_MAC_37_15);
	MAC_38_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_0, data_out=>output_MAC_38_0);
	MAC_38_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_1, data_out=>output_MAC_38_1);
	MAC_38_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_2, data_out=>output_MAC_38_2);
	MAC_38_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_3, data_out=>output_MAC_38_3);
	MAC_38_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_4, data_out=>output_MAC_38_4);
	MAC_38_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_5, data_out=>output_MAC_38_5);
	MAC_38_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_6, data_out=>output_MAC_38_6);
	MAC_38_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_7, data_out=>output_MAC_38_7);
	MAC_38_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_8, data_out=>output_MAC_38_8);
	MAC_38_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_9, data_out=>output_MAC_38_9);
	MAC_38_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_10, data_out=>output_MAC_38_10);
	MAC_38_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_11, data_out=>output_MAC_38_11);
	MAC_38_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_12, data_out=>output_MAC_38_12);
	MAC_38_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_13, data_out=>output_MAC_38_13);
	MAC_38_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_14, data_out=>output_MAC_38_14);
	MAC_38_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_38, data_in_B=>input_col_15, data_out=>output_MAC_38_15);
	MAC_39_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_0, data_out=>output_MAC_39_0);
	MAC_39_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_1, data_out=>output_MAC_39_1);
	MAC_39_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_2, data_out=>output_MAC_39_2);
	MAC_39_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_3, data_out=>output_MAC_39_3);
	MAC_39_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_4, data_out=>output_MAC_39_4);
	MAC_39_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_5, data_out=>output_MAC_39_5);
	MAC_39_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_6, data_out=>output_MAC_39_6);
	MAC_39_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_7, data_out=>output_MAC_39_7);
	MAC_39_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_8, data_out=>output_MAC_39_8);
	MAC_39_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_9, data_out=>output_MAC_39_9);
	MAC_39_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_10, data_out=>output_MAC_39_10);
	MAC_39_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_11, data_out=>output_MAC_39_11);
	MAC_39_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_12, data_out=>output_MAC_39_12);
	MAC_39_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_13, data_out=>output_MAC_39_13);
	MAC_39_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_14, data_out=>output_MAC_39_14);
	MAC_39_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_39, data_in_B=>input_col_15, data_out=>output_MAC_39_15);
	MAC_40_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_0, data_out=>output_MAC_40_0);
	MAC_40_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_1, data_out=>output_MAC_40_1);
	MAC_40_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_2, data_out=>output_MAC_40_2);
	MAC_40_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_3, data_out=>output_MAC_40_3);
	MAC_40_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_4, data_out=>output_MAC_40_4);
	MAC_40_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_5, data_out=>output_MAC_40_5);
	MAC_40_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_6, data_out=>output_MAC_40_6);
	MAC_40_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_7, data_out=>output_MAC_40_7);
	MAC_40_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_8, data_out=>output_MAC_40_8);
	MAC_40_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_9, data_out=>output_MAC_40_9);
	MAC_40_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_10, data_out=>output_MAC_40_10);
	MAC_40_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_11, data_out=>output_MAC_40_11);
	MAC_40_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_12, data_out=>output_MAC_40_12);
	MAC_40_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_13, data_out=>output_MAC_40_13);
	MAC_40_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_14, data_out=>output_MAC_40_14);
	MAC_40_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_40, data_in_B=>input_col_15, data_out=>output_MAC_40_15);
	MAC_41_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_0, data_out=>output_MAC_41_0);
	MAC_41_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_1, data_out=>output_MAC_41_1);
	MAC_41_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_2, data_out=>output_MAC_41_2);
	MAC_41_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_3, data_out=>output_MAC_41_3);
	MAC_41_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_4, data_out=>output_MAC_41_4);
	MAC_41_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_5, data_out=>output_MAC_41_5);
	MAC_41_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_6, data_out=>output_MAC_41_6);
	MAC_41_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_7, data_out=>output_MAC_41_7);
	MAC_41_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_8, data_out=>output_MAC_41_8);
	MAC_41_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_9, data_out=>output_MAC_41_9);
	MAC_41_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_10, data_out=>output_MAC_41_10);
	MAC_41_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_11, data_out=>output_MAC_41_11);
	MAC_41_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_12, data_out=>output_MAC_41_12);
	MAC_41_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_13, data_out=>output_MAC_41_13);
	MAC_41_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_14, data_out=>output_MAC_41_14);
	MAC_41_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_41, data_in_B=>input_col_15, data_out=>output_MAC_41_15);
	MAC_42_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_0, data_out=>output_MAC_42_0);
	MAC_42_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_1, data_out=>output_MAC_42_1);
	MAC_42_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_2, data_out=>output_MAC_42_2);
	MAC_42_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_3, data_out=>output_MAC_42_3);
	MAC_42_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_4, data_out=>output_MAC_42_4);
	MAC_42_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_5, data_out=>output_MAC_42_5);
	MAC_42_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_6, data_out=>output_MAC_42_6);
	MAC_42_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_7, data_out=>output_MAC_42_7);
	MAC_42_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_8, data_out=>output_MAC_42_8);
	MAC_42_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_9, data_out=>output_MAC_42_9);
	MAC_42_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_10, data_out=>output_MAC_42_10);
	MAC_42_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_11, data_out=>output_MAC_42_11);
	MAC_42_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_12, data_out=>output_MAC_42_12);
	MAC_42_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_13, data_out=>output_MAC_42_13);
	MAC_42_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_14, data_out=>output_MAC_42_14);
	MAC_42_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_42, data_in_B=>input_col_15, data_out=>output_MAC_42_15);
	MAC_43_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_0, data_out=>output_MAC_43_0);
	MAC_43_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_1, data_out=>output_MAC_43_1);
	MAC_43_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_2, data_out=>output_MAC_43_2);
	MAC_43_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_3, data_out=>output_MAC_43_3);
	MAC_43_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_4, data_out=>output_MAC_43_4);
	MAC_43_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_5, data_out=>output_MAC_43_5);
	MAC_43_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_6, data_out=>output_MAC_43_6);
	MAC_43_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_7, data_out=>output_MAC_43_7);
	MAC_43_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_8, data_out=>output_MAC_43_8);
	MAC_43_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_9, data_out=>output_MAC_43_9);
	MAC_43_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_10, data_out=>output_MAC_43_10);
	MAC_43_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_11, data_out=>output_MAC_43_11);
	MAC_43_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_12, data_out=>output_MAC_43_12);
	MAC_43_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_13, data_out=>output_MAC_43_13);
	MAC_43_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_14, data_out=>output_MAC_43_14);
	MAC_43_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_43, data_in_B=>input_col_15, data_out=>output_MAC_43_15);
	MAC_44_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_0, data_out=>output_MAC_44_0);
	MAC_44_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_1, data_out=>output_MAC_44_1);
	MAC_44_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_2, data_out=>output_MAC_44_2);
	MAC_44_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_3, data_out=>output_MAC_44_3);
	MAC_44_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_4, data_out=>output_MAC_44_4);
	MAC_44_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_5, data_out=>output_MAC_44_5);
	MAC_44_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_6, data_out=>output_MAC_44_6);
	MAC_44_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_7, data_out=>output_MAC_44_7);
	MAC_44_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_8, data_out=>output_MAC_44_8);
	MAC_44_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_9, data_out=>output_MAC_44_9);
	MAC_44_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_10, data_out=>output_MAC_44_10);
	MAC_44_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_11, data_out=>output_MAC_44_11);
	MAC_44_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_12, data_out=>output_MAC_44_12);
	MAC_44_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_13, data_out=>output_MAC_44_13);
	MAC_44_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_14, data_out=>output_MAC_44_14);
	MAC_44_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_44, data_in_B=>input_col_15, data_out=>output_MAC_44_15);
	MAC_45_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_0, data_out=>output_MAC_45_0);
	MAC_45_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_1, data_out=>output_MAC_45_1);
	MAC_45_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_2, data_out=>output_MAC_45_2);
	MAC_45_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_3, data_out=>output_MAC_45_3);
	MAC_45_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_4, data_out=>output_MAC_45_4);
	MAC_45_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_5, data_out=>output_MAC_45_5);
	MAC_45_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_6, data_out=>output_MAC_45_6);
	MAC_45_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_7, data_out=>output_MAC_45_7);
	MAC_45_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_8, data_out=>output_MAC_45_8);
	MAC_45_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_9, data_out=>output_MAC_45_9);
	MAC_45_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_10, data_out=>output_MAC_45_10);
	MAC_45_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_11, data_out=>output_MAC_45_11);
	MAC_45_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_12, data_out=>output_MAC_45_12);
	MAC_45_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_13, data_out=>output_MAC_45_13);
	MAC_45_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_14, data_out=>output_MAC_45_14);
	MAC_45_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_45, data_in_B=>input_col_15, data_out=>output_MAC_45_15);
	MAC_46_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_0, data_out=>output_MAC_46_0);
	MAC_46_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_1, data_out=>output_MAC_46_1);
	MAC_46_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_2, data_out=>output_MAC_46_2);
	MAC_46_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_3, data_out=>output_MAC_46_3);
	MAC_46_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_4, data_out=>output_MAC_46_4);
	MAC_46_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_5, data_out=>output_MAC_46_5);
	MAC_46_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_6, data_out=>output_MAC_46_6);
	MAC_46_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_7, data_out=>output_MAC_46_7);
	MAC_46_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_8, data_out=>output_MAC_46_8);
	MAC_46_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_9, data_out=>output_MAC_46_9);
	MAC_46_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_10, data_out=>output_MAC_46_10);
	MAC_46_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_11, data_out=>output_MAC_46_11);
	MAC_46_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_12, data_out=>output_MAC_46_12);
	MAC_46_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_13, data_out=>output_MAC_46_13);
	MAC_46_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_14, data_out=>output_MAC_46_14);
	MAC_46_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_46, data_in_B=>input_col_15, data_out=>output_MAC_46_15);
	MAC_47_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_0, data_out=>output_MAC_47_0);
	MAC_47_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_1, data_out=>output_MAC_47_1);
	MAC_47_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_2, data_out=>output_MAC_47_2);
	MAC_47_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_3, data_out=>output_MAC_47_3);
	MAC_47_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_4, data_out=>output_MAC_47_4);
	MAC_47_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_5, data_out=>output_MAC_47_5);
	MAC_47_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_6, data_out=>output_MAC_47_6);
	MAC_47_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_7, data_out=>output_MAC_47_7);
	MAC_47_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_8, data_out=>output_MAC_47_8);
	MAC_47_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_9, data_out=>output_MAC_47_9);
	MAC_47_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_10, data_out=>output_MAC_47_10);
	MAC_47_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_11, data_out=>output_MAC_47_11);
	MAC_47_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_12, data_out=>output_MAC_47_12);
	MAC_47_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_13, data_out=>output_MAC_47_13);
	MAC_47_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_14, data_out=>output_MAC_47_14);
	MAC_47_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_47, data_in_B=>input_col_15, data_out=>output_MAC_47_15);
	MAC_48_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_0, data_out=>output_MAC_48_0);
	MAC_48_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_1, data_out=>output_MAC_48_1);
	MAC_48_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_2, data_out=>output_MAC_48_2);
	MAC_48_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_3, data_out=>output_MAC_48_3);
	MAC_48_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_4, data_out=>output_MAC_48_4);
	MAC_48_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_5, data_out=>output_MAC_48_5);
	MAC_48_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_6, data_out=>output_MAC_48_6);
	MAC_48_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_7, data_out=>output_MAC_48_7);
	MAC_48_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_8, data_out=>output_MAC_48_8);
	MAC_48_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_9, data_out=>output_MAC_48_9);
	MAC_48_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_10, data_out=>output_MAC_48_10);
	MAC_48_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_11, data_out=>output_MAC_48_11);
	MAC_48_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_12, data_out=>output_MAC_48_12);
	MAC_48_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_13, data_out=>output_MAC_48_13);
	MAC_48_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_14, data_out=>output_MAC_48_14);
	MAC_48_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_48, data_in_B=>input_col_15, data_out=>output_MAC_48_15);
	MAC_49_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_0, data_out=>output_MAC_49_0);
	MAC_49_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_1, data_out=>output_MAC_49_1);
	MAC_49_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_2, data_out=>output_MAC_49_2);
	MAC_49_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_3, data_out=>output_MAC_49_3);
	MAC_49_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_4, data_out=>output_MAC_49_4);
	MAC_49_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_5, data_out=>output_MAC_49_5);
	MAC_49_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_6, data_out=>output_MAC_49_6);
	MAC_49_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_7, data_out=>output_MAC_49_7);
	MAC_49_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_8, data_out=>output_MAC_49_8);
	MAC_49_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_9, data_out=>output_MAC_49_9);
	MAC_49_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_10, data_out=>output_MAC_49_10);
	MAC_49_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_11, data_out=>output_MAC_49_11);
	MAC_49_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_12, data_out=>output_MAC_49_12);
	MAC_49_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_13, data_out=>output_MAC_49_13);
	MAC_49_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_14, data_out=>output_MAC_49_14);
	MAC_49_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_49, data_in_B=>input_col_15, data_out=>output_MAC_49_15);
	MAC_50_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_0, data_out=>output_MAC_50_0);
	MAC_50_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_1, data_out=>output_MAC_50_1);
	MAC_50_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_2, data_out=>output_MAC_50_2);
	MAC_50_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_3, data_out=>output_MAC_50_3);
	MAC_50_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_4, data_out=>output_MAC_50_4);
	MAC_50_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_5, data_out=>output_MAC_50_5);
	MAC_50_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_6, data_out=>output_MAC_50_6);
	MAC_50_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_7, data_out=>output_MAC_50_7);
	MAC_50_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_8, data_out=>output_MAC_50_8);
	MAC_50_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_9, data_out=>output_MAC_50_9);
	MAC_50_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_10, data_out=>output_MAC_50_10);
	MAC_50_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_11, data_out=>output_MAC_50_11);
	MAC_50_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_12, data_out=>output_MAC_50_12);
	MAC_50_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_13, data_out=>output_MAC_50_13);
	MAC_50_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_14, data_out=>output_MAC_50_14);
	MAC_50_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_50, data_in_B=>input_col_15, data_out=>output_MAC_50_15);
	MAC_51_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_0, data_out=>output_MAC_51_0);
	MAC_51_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_1, data_out=>output_MAC_51_1);
	MAC_51_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_2, data_out=>output_MAC_51_2);
	MAC_51_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_3, data_out=>output_MAC_51_3);
	MAC_51_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_4, data_out=>output_MAC_51_4);
	MAC_51_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_5, data_out=>output_MAC_51_5);
	MAC_51_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_6, data_out=>output_MAC_51_6);
	MAC_51_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_7, data_out=>output_MAC_51_7);
	MAC_51_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_8, data_out=>output_MAC_51_8);
	MAC_51_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_9, data_out=>output_MAC_51_9);
	MAC_51_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_10, data_out=>output_MAC_51_10);
	MAC_51_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_11, data_out=>output_MAC_51_11);
	MAC_51_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_12, data_out=>output_MAC_51_12);
	MAC_51_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_13, data_out=>output_MAC_51_13);
	MAC_51_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_14, data_out=>output_MAC_51_14);
	MAC_51_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_51, data_in_B=>input_col_15, data_out=>output_MAC_51_15);
	MAC_52_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_0, data_out=>output_MAC_52_0);
	MAC_52_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_1, data_out=>output_MAC_52_1);
	MAC_52_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_2, data_out=>output_MAC_52_2);
	MAC_52_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_3, data_out=>output_MAC_52_3);
	MAC_52_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_4, data_out=>output_MAC_52_4);
	MAC_52_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_5, data_out=>output_MAC_52_5);
	MAC_52_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_6, data_out=>output_MAC_52_6);
	MAC_52_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_7, data_out=>output_MAC_52_7);
	MAC_52_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_8, data_out=>output_MAC_52_8);
	MAC_52_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_9, data_out=>output_MAC_52_9);
	MAC_52_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_10, data_out=>output_MAC_52_10);
	MAC_52_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_11, data_out=>output_MAC_52_11);
	MAC_52_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_12, data_out=>output_MAC_52_12);
	MAC_52_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_13, data_out=>output_MAC_52_13);
	MAC_52_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_14, data_out=>output_MAC_52_14);
	MAC_52_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_52, data_in_B=>input_col_15, data_out=>output_MAC_52_15);
	MAC_53_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_0, data_out=>output_MAC_53_0);
	MAC_53_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_1, data_out=>output_MAC_53_1);
	MAC_53_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_2, data_out=>output_MAC_53_2);
	MAC_53_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_3, data_out=>output_MAC_53_3);
	MAC_53_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_4, data_out=>output_MAC_53_4);
	MAC_53_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_5, data_out=>output_MAC_53_5);
	MAC_53_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_6, data_out=>output_MAC_53_6);
	MAC_53_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_7, data_out=>output_MAC_53_7);
	MAC_53_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_8, data_out=>output_MAC_53_8);
	MAC_53_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_9, data_out=>output_MAC_53_9);
	MAC_53_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_10, data_out=>output_MAC_53_10);
	MAC_53_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_11, data_out=>output_MAC_53_11);
	MAC_53_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_12, data_out=>output_MAC_53_12);
	MAC_53_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_13, data_out=>output_MAC_53_13);
	MAC_53_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_14, data_out=>output_MAC_53_14);
	MAC_53_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_53, data_in_B=>input_col_15, data_out=>output_MAC_53_15);
	MAC_54_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_0, data_out=>output_MAC_54_0);
	MAC_54_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_1, data_out=>output_MAC_54_1);
	MAC_54_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_2, data_out=>output_MAC_54_2);
	MAC_54_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_3, data_out=>output_MAC_54_3);
	MAC_54_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_4, data_out=>output_MAC_54_4);
	MAC_54_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_5, data_out=>output_MAC_54_5);
	MAC_54_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_6, data_out=>output_MAC_54_6);
	MAC_54_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_7, data_out=>output_MAC_54_7);
	MAC_54_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_8, data_out=>output_MAC_54_8);
	MAC_54_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_9, data_out=>output_MAC_54_9);
	MAC_54_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_10, data_out=>output_MAC_54_10);
	MAC_54_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_11, data_out=>output_MAC_54_11);
	MAC_54_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_12, data_out=>output_MAC_54_12);
	MAC_54_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_13, data_out=>output_MAC_54_13);
	MAC_54_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_14, data_out=>output_MAC_54_14);
	MAC_54_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_54, data_in_B=>input_col_15, data_out=>output_MAC_54_15);
	MAC_55_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_0, data_out=>output_MAC_55_0);
	MAC_55_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_1, data_out=>output_MAC_55_1);
	MAC_55_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_2, data_out=>output_MAC_55_2);
	MAC_55_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_3, data_out=>output_MAC_55_3);
	MAC_55_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_4, data_out=>output_MAC_55_4);
	MAC_55_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_5, data_out=>output_MAC_55_5);
	MAC_55_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_6, data_out=>output_MAC_55_6);
	MAC_55_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_7, data_out=>output_MAC_55_7);
	MAC_55_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_8, data_out=>output_MAC_55_8);
	MAC_55_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_9, data_out=>output_MAC_55_9);
	MAC_55_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_10, data_out=>output_MAC_55_10);
	MAC_55_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_11, data_out=>output_MAC_55_11);
	MAC_55_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_12, data_out=>output_MAC_55_12);
	MAC_55_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_13, data_out=>output_MAC_55_13);
	MAC_55_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_14, data_out=>output_MAC_55_14);
	MAC_55_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_55, data_in_B=>input_col_15, data_out=>output_MAC_55_15);
	MAC_56_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_0, data_out=>output_MAC_56_0);
	MAC_56_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_1, data_out=>output_MAC_56_1);
	MAC_56_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_2, data_out=>output_MAC_56_2);
	MAC_56_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_3, data_out=>output_MAC_56_3);
	MAC_56_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_4, data_out=>output_MAC_56_4);
	MAC_56_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_5, data_out=>output_MAC_56_5);
	MAC_56_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_6, data_out=>output_MAC_56_6);
	MAC_56_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_7, data_out=>output_MAC_56_7);
	MAC_56_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_8, data_out=>output_MAC_56_8);
	MAC_56_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_9, data_out=>output_MAC_56_9);
	MAC_56_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_10, data_out=>output_MAC_56_10);
	MAC_56_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_11, data_out=>output_MAC_56_11);
	MAC_56_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_12, data_out=>output_MAC_56_12);
	MAC_56_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_13, data_out=>output_MAC_56_13);
	MAC_56_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_14, data_out=>output_MAC_56_14);
	MAC_56_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_56, data_in_B=>input_col_15, data_out=>output_MAC_56_15);
	MAC_57_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_0, data_out=>output_MAC_57_0);
	MAC_57_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_1, data_out=>output_MAC_57_1);
	MAC_57_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_2, data_out=>output_MAC_57_2);
	MAC_57_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_3, data_out=>output_MAC_57_3);
	MAC_57_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_4, data_out=>output_MAC_57_4);
	MAC_57_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_5, data_out=>output_MAC_57_5);
	MAC_57_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_6, data_out=>output_MAC_57_6);
	MAC_57_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_7, data_out=>output_MAC_57_7);
	MAC_57_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_8, data_out=>output_MAC_57_8);
	MAC_57_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_9, data_out=>output_MAC_57_9);
	MAC_57_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_10, data_out=>output_MAC_57_10);
	MAC_57_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_11, data_out=>output_MAC_57_11);
	MAC_57_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_12, data_out=>output_MAC_57_12);
	MAC_57_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_13, data_out=>output_MAC_57_13);
	MAC_57_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_14, data_out=>output_MAC_57_14);
	MAC_57_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_57, data_in_B=>input_col_15, data_out=>output_MAC_57_15);
	MAC_58_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_0, data_out=>output_MAC_58_0);
	MAC_58_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_1, data_out=>output_MAC_58_1);
	MAC_58_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_2, data_out=>output_MAC_58_2);
	MAC_58_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_3, data_out=>output_MAC_58_3);
	MAC_58_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_4, data_out=>output_MAC_58_4);
	MAC_58_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_5, data_out=>output_MAC_58_5);
	MAC_58_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_6, data_out=>output_MAC_58_6);
	MAC_58_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_7, data_out=>output_MAC_58_7);
	MAC_58_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_8, data_out=>output_MAC_58_8);
	MAC_58_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_9, data_out=>output_MAC_58_9);
	MAC_58_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_10, data_out=>output_MAC_58_10);
	MAC_58_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_11, data_out=>output_MAC_58_11);
	MAC_58_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_12, data_out=>output_MAC_58_12);
	MAC_58_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_13, data_out=>output_MAC_58_13);
	MAC_58_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_14, data_out=>output_MAC_58_14);
	MAC_58_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_58, data_in_B=>input_col_15, data_out=>output_MAC_58_15);
	MAC_59_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_0, data_out=>output_MAC_59_0);
	MAC_59_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_1, data_out=>output_MAC_59_1);
	MAC_59_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_2, data_out=>output_MAC_59_2);
	MAC_59_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_3, data_out=>output_MAC_59_3);
	MAC_59_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_4, data_out=>output_MAC_59_4);
	MAC_59_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_5, data_out=>output_MAC_59_5);
	MAC_59_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_6, data_out=>output_MAC_59_6);
	MAC_59_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_7, data_out=>output_MAC_59_7);
	MAC_59_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_8, data_out=>output_MAC_59_8);
	MAC_59_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_9, data_out=>output_MAC_59_9);
	MAC_59_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_10, data_out=>output_MAC_59_10);
	MAC_59_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_11, data_out=>output_MAC_59_11);
	MAC_59_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_12, data_out=>output_MAC_59_12);
	MAC_59_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_13, data_out=>output_MAC_59_13);
	MAC_59_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_14, data_out=>output_MAC_59_14);
	MAC_59_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_59, data_in_B=>input_col_15, data_out=>output_MAC_59_15);
	MAC_60_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_0, data_out=>output_MAC_60_0);
	MAC_60_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_1, data_out=>output_MAC_60_1);
	MAC_60_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_2, data_out=>output_MAC_60_2);
	MAC_60_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_3, data_out=>output_MAC_60_3);
	MAC_60_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_4, data_out=>output_MAC_60_4);
	MAC_60_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_5, data_out=>output_MAC_60_5);
	MAC_60_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_6, data_out=>output_MAC_60_6);
	MAC_60_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_7, data_out=>output_MAC_60_7);
	MAC_60_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_8, data_out=>output_MAC_60_8);
	MAC_60_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_9, data_out=>output_MAC_60_9);
	MAC_60_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_10, data_out=>output_MAC_60_10);
	MAC_60_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_11, data_out=>output_MAC_60_11);
	MAC_60_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_12, data_out=>output_MAC_60_12);
	MAC_60_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_13, data_out=>output_MAC_60_13);
	MAC_60_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_14, data_out=>output_MAC_60_14);
	MAC_60_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_60, data_in_B=>input_col_15, data_out=>output_MAC_60_15);
	MAC_61_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_0, data_out=>output_MAC_61_0);
	MAC_61_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_1, data_out=>output_MAC_61_1);
	MAC_61_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_2, data_out=>output_MAC_61_2);
	MAC_61_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_3, data_out=>output_MAC_61_3);
	MAC_61_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_4, data_out=>output_MAC_61_4);
	MAC_61_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_5, data_out=>output_MAC_61_5);
	MAC_61_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_6, data_out=>output_MAC_61_6);
	MAC_61_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_7, data_out=>output_MAC_61_7);
	MAC_61_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_8, data_out=>output_MAC_61_8);
	MAC_61_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_9, data_out=>output_MAC_61_9);
	MAC_61_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_10, data_out=>output_MAC_61_10);
	MAC_61_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_11, data_out=>output_MAC_61_11);
	MAC_61_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_12, data_out=>output_MAC_61_12);
	MAC_61_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_13, data_out=>output_MAC_61_13);
	MAC_61_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_14, data_out=>output_MAC_61_14);
	MAC_61_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_61, data_in_B=>input_col_15, data_out=>output_MAC_61_15);
	MAC_62_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_0, data_out=>output_MAC_62_0);
	MAC_62_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_1, data_out=>output_MAC_62_1);
	MAC_62_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_2, data_out=>output_MAC_62_2);
	MAC_62_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_3, data_out=>output_MAC_62_3);
	MAC_62_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_4, data_out=>output_MAC_62_4);
	MAC_62_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_5, data_out=>output_MAC_62_5);
	MAC_62_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_6, data_out=>output_MAC_62_6);
	MAC_62_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_7, data_out=>output_MAC_62_7);
	MAC_62_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_8, data_out=>output_MAC_62_8);
	MAC_62_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_9, data_out=>output_MAC_62_9);
	MAC_62_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_10, data_out=>output_MAC_62_10);
	MAC_62_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_11, data_out=>output_MAC_62_11);
	MAC_62_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_12, data_out=>output_MAC_62_12);
	MAC_62_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_13, data_out=>output_MAC_62_13);
	MAC_62_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_14, data_out=>output_MAC_62_14);
	MAC_62_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_62, data_in_B=>input_col_15, data_out=>output_MAC_62_15);
	MAC_63_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_0, data_out=>output_MAC_63_0);
	MAC_63_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_1, data_out=>output_MAC_63_1);
	MAC_63_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_2, data_out=>output_MAC_63_2);
	MAC_63_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_3, data_out=>output_MAC_63_3);
	MAC_63_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_4, data_out=>output_MAC_63_4);
	MAC_63_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_5, data_out=>output_MAC_63_5);
	MAC_63_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_6, data_out=>output_MAC_63_6);
	MAC_63_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_7, data_out=>output_MAC_63_7);
	MAC_63_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_8, data_out=>output_MAC_63_8);
	MAC_63_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_9, data_out=>output_MAC_63_9);
	MAC_63_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_10, data_out=>output_MAC_63_10);
	MAC_63_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_11, data_out=>output_MAC_63_11);
	MAC_63_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_12, data_out=>output_MAC_63_12);
	MAC_63_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_13, data_out=>output_MAC_63_13);
	MAC_63_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_14, data_out=>output_MAC_63_14);
	MAC_63_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_63, data_in_B=>input_col_15, data_out=>output_MAC_63_15);

	mux_row_0: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_0_0, I1=>output_MAC_0_1, I2=>output_MAC_0_2, I3=>output_MAC_0_3, I4=>output_MAC_0_4, I5=>output_MAC_0_5, I6=>output_MAC_0_6, I7=>output_MAC_0_7, I8=>output_MAC_0_8, I9=>output_MAC_0_9, I10=>output_MAC_0_10, I11=>output_MAC_0_11, I12=>output_MAC_0_12, I13=>output_MAC_0_13, I14=>output_MAC_0_14, I15=>output_MAC_0_15, 
		SEL_mux=>SEL_mux, O=>output_row_0);

	mux_row_1: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_1_0, I1=>output_MAC_1_1, I2=>output_MAC_1_2, I3=>output_MAC_1_3, I4=>output_MAC_1_4, I5=>output_MAC_1_5, I6=>output_MAC_1_6, I7=>output_MAC_1_7, I8=>output_MAC_1_8, I9=>output_MAC_1_9, I10=>output_MAC_1_10, I11=>output_MAC_1_11, I12=>output_MAC_1_12, I13=>output_MAC_1_13, I14=>output_MAC_1_14, I15=>output_MAC_1_15, 
		SEL_mux=>SEL_mux, O=>output_row_1);

	mux_row_2: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_2_0, I1=>output_MAC_2_1, I2=>output_MAC_2_2, I3=>output_MAC_2_3, I4=>output_MAC_2_4, I5=>output_MAC_2_5, I6=>output_MAC_2_6, I7=>output_MAC_2_7, I8=>output_MAC_2_8, I9=>output_MAC_2_9, I10=>output_MAC_2_10, I11=>output_MAC_2_11, I12=>output_MAC_2_12, I13=>output_MAC_2_13, I14=>output_MAC_2_14, I15=>output_MAC_2_15, 
		SEL_mux=>SEL_mux, O=>output_row_2);

	mux_row_3: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_3_0, I1=>output_MAC_3_1, I2=>output_MAC_3_2, I3=>output_MAC_3_3, I4=>output_MAC_3_4, I5=>output_MAC_3_5, I6=>output_MAC_3_6, I7=>output_MAC_3_7, I8=>output_MAC_3_8, I9=>output_MAC_3_9, I10=>output_MAC_3_10, I11=>output_MAC_3_11, I12=>output_MAC_3_12, I13=>output_MAC_3_13, I14=>output_MAC_3_14, I15=>output_MAC_3_15, 
		SEL_mux=>SEL_mux, O=>output_row_3);

	mux_row_4: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_4_0, I1=>output_MAC_4_1, I2=>output_MAC_4_2, I3=>output_MAC_4_3, I4=>output_MAC_4_4, I5=>output_MAC_4_5, I6=>output_MAC_4_6, I7=>output_MAC_4_7, I8=>output_MAC_4_8, I9=>output_MAC_4_9, I10=>output_MAC_4_10, I11=>output_MAC_4_11, I12=>output_MAC_4_12, I13=>output_MAC_4_13, I14=>output_MAC_4_14, I15=>output_MAC_4_15, 
		SEL_mux=>SEL_mux, O=>output_row_4);

	mux_row_5: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_5_0, I1=>output_MAC_5_1, I2=>output_MAC_5_2, I3=>output_MAC_5_3, I4=>output_MAC_5_4, I5=>output_MAC_5_5, I6=>output_MAC_5_6, I7=>output_MAC_5_7, I8=>output_MAC_5_8, I9=>output_MAC_5_9, I10=>output_MAC_5_10, I11=>output_MAC_5_11, I12=>output_MAC_5_12, I13=>output_MAC_5_13, I14=>output_MAC_5_14, I15=>output_MAC_5_15, 
		SEL_mux=>SEL_mux, O=>output_row_5);

	mux_row_6: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_6_0, I1=>output_MAC_6_1, I2=>output_MAC_6_2, I3=>output_MAC_6_3, I4=>output_MAC_6_4, I5=>output_MAC_6_5, I6=>output_MAC_6_6, I7=>output_MAC_6_7, I8=>output_MAC_6_8, I9=>output_MAC_6_9, I10=>output_MAC_6_10, I11=>output_MAC_6_11, I12=>output_MAC_6_12, I13=>output_MAC_6_13, I14=>output_MAC_6_14, I15=>output_MAC_6_15, 
		SEL_mux=>SEL_mux, O=>output_row_6);

	mux_row_7: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_7_0, I1=>output_MAC_7_1, I2=>output_MAC_7_2, I3=>output_MAC_7_3, I4=>output_MAC_7_4, I5=>output_MAC_7_5, I6=>output_MAC_7_6, I7=>output_MAC_7_7, I8=>output_MAC_7_8, I9=>output_MAC_7_9, I10=>output_MAC_7_10, I11=>output_MAC_7_11, I12=>output_MAC_7_12, I13=>output_MAC_7_13, I14=>output_MAC_7_14, I15=>output_MAC_7_15, 
		SEL_mux=>SEL_mux, O=>output_row_7);

	mux_row_8: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_8_0, I1=>output_MAC_8_1, I2=>output_MAC_8_2, I3=>output_MAC_8_3, I4=>output_MAC_8_4, I5=>output_MAC_8_5, I6=>output_MAC_8_6, I7=>output_MAC_8_7, I8=>output_MAC_8_8, I9=>output_MAC_8_9, I10=>output_MAC_8_10, I11=>output_MAC_8_11, I12=>output_MAC_8_12, I13=>output_MAC_8_13, I14=>output_MAC_8_14, I15=>output_MAC_8_15, 
		SEL_mux=>SEL_mux, O=>output_row_8);

	mux_row_9: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_9_0, I1=>output_MAC_9_1, I2=>output_MAC_9_2, I3=>output_MAC_9_3, I4=>output_MAC_9_4, I5=>output_MAC_9_5, I6=>output_MAC_9_6, I7=>output_MAC_9_7, I8=>output_MAC_9_8, I9=>output_MAC_9_9, I10=>output_MAC_9_10, I11=>output_MAC_9_11, I12=>output_MAC_9_12, I13=>output_MAC_9_13, I14=>output_MAC_9_14, I15=>output_MAC_9_15, 
		SEL_mux=>SEL_mux, O=>output_row_9);

	mux_row_10: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_10_0, I1=>output_MAC_10_1, I2=>output_MAC_10_2, I3=>output_MAC_10_3, I4=>output_MAC_10_4, I5=>output_MAC_10_5, I6=>output_MAC_10_6, I7=>output_MAC_10_7, I8=>output_MAC_10_8, I9=>output_MAC_10_9, I10=>output_MAC_10_10, I11=>output_MAC_10_11, I12=>output_MAC_10_12, I13=>output_MAC_10_13, I14=>output_MAC_10_14, I15=>output_MAC_10_15, 
		SEL_mux=>SEL_mux, O=>output_row_10);

	mux_row_11: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_11_0, I1=>output_MAC_11_1, I2=>output_MAC_11_2, I3=>output_MAC_11_3, I4=>output_MAC_11_4, I5=>output_MAC_11_5, I6=>output_MAC_11_6, I7=>output_MAC_11_7, I8=>output_MAC_11_8, I9=>output_MAC_11_9, I10=>output_MAC_11_10, I11=>output_MAC_11_11, I12=>output_MAC_11_12, I13=>output_MAC_11_13, I14=>output_MAC_11_14, I15=>output_MAC_11_15, 
		SEL_mux=>SEL_mux, O=>output_row_11);

	mux_row_12: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_12_0, I1=>output_MAC_12_1, I2=>output_MAC_12_2, I3=>output_MAC_12_3, I4=>output_MAC_12_4, I5=>output_MAC_12_5, I6=>output_MAC_12_6, I7=>output_MAC_12_7, I8=>output_MAC_12_8, I9=>output_MAC_12_9, I10=>output_MAC_12_10, I11=>output_MAC_12_11, I12=>output_MAC_12_12, I13=>output_MAC_12_13, I14=>output_MAC_12_14, I15=>output_MAC_12_15, 
		SEL_mux=>SEL_mux, O=>output_row_12);

	mux_row_13: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_13_0, I1=>output_MAC_13_1, I2=>output_MAC_13_2, I3=>output_MAC_13_3, I4=>output_MAC_13_4, I5=>output_MAC_13_5, I6=>output_MAC_13_6, I7=>output_MAC_13_7, I8=>output_MAC_13_8, I9=>output_MAC_13_9, I10=>output_MAC_13_10, I11=>output_MAC_13_11, I12=>output_MAC_13_12, I13=>output_MAC_13_13, I14=>output_MAC_13_14, I15=>output_MAC_13_15, 
		SEL_mux=>SEL_mux, O=>output_row_13);

	mux_row_14: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_14_0, I1=>output_MAC_14_1, I2=>output_MAC_14_2, I3=>output_MAC_14_3, I4=>output_MAC_14_4, I5=>output_MAC_14_5, I6=>output_MAC_14_6, I7=>output_MAC_14_7, I8=>output_MAC_14_8, I9=>output_MAC_14_9, I10=>output_MAC_14_10, I11=>output_MAC_14_11, I12=>output_MAC_14_12, I13=>output_MAC_14_13, I14=>output_MAC_14_14, I15=>output_MAC_14_15, 
		SEL_mux=>SEL_mux, O=>output_row_14);

	mux_row_15: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_15_0, I1=>output_MAC_15_1, I2=>output_MAC_15_2, I3=>output_MAC_15_3, I4=>output_MAC_15_4, I5=>output_MAC_15_5, I6=>output_MAC_15_6, I7=>output_MAC_15_7, I8=>output_MAC_15_8, I9=>output_MAC_15_9, I10=>output_MAC_15_10, I11=>output_MAC_15_11, I12=>output_MAC_15_12, I13=>output_MAC_15_13, I14=>output_MAC_15_14, I15=>output_MAC_15_15, 
		SEL_mux=>SEL_mux, O=>output_row_15);

	mux_row_16: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_16_0, I1=>output_MAC_16_1, I2=>output_MAC_16_2, I3=>output_MAC_16_3, I4=>output_MAC_16_4, I5=>output_MAC_16_5, I6=>output_MAC_16_6, I7=>output_MAC_16_7, I8=>output_MAC_16_8, I9=>output_MAC_16_9, I10=>output_MAC_16_10, I11=>output_MAC_16_11, I12=>output_MAC_16_12, I13=>output_MAC_16_13, I14=>output_MAC_16_14, I15=>output_MAC_16_15, 
		SEL_mux=>SEL_mux, O=>output_row_16);

	mux_row_17: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_17_0, I1=>output_MAC_17_1, I2=>output_MAC_17_2, I3=>output_MAC_17_3, I4=>output_MAC_17_4, I5=>output_MAC_17_5, I6=>output_MAC_17_6, I7=>output_MAC_17_7, I8=>output_MAC_17_8, I9=>output_MAC_17_9, I10=>output_MAC_17_10, I11=>output_MAC_17_11, I12=>output_MAC_17_12, I13=>output_MAC_17_13, I14=>output_MAC_17_14, I15=>output_MAC_17_15, 
		SEL_mux=>SEL_mux, O=>output_row_17);

	mux_row_18: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_18_0, I1=>output_MAC_18_1, I2=>output_MAC_18_2, I3=>output_MAC_18_3, I4=>output_MAC_18_4, I5=>output_MAC_18_5, I6=>output_MAC_18_6, I7=>output_MAC_18_7, I8=>output_MAC_18_8, I9=>output_MAC_18_9, I10=>output_MAC_18_10, I11=>output_MAC_18_11, I12=>output_MAC_18_12, I13=>output_MAC_18_13, I14=>output_MAC_18_14, I15=>output_MAC_18_15, 
		SEL_mux=>SEL_mux, O=>output_row_18);

	mux_row_19: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_19_0, I1=>output_MAC_19_1, I2=>output_MAC_19_2, I3=>output_MAC_19_3, I4=>output_MAC_19_4, I5=>output_MAC_19_5, I6=>output_MAC_19_6, I7=>output_MAC_19_7, I8=>output_MAC_19_8, I9=>output_MAC_19_9, I10=>output_MAC_19_10, I11=>output_MAC_19_11, I12=>output_MAC_19_12, I13=>output_MAC_19_13, I14=>output_MAC_19_14, I15=>output_MAC_19_15, 
		SEL_mux=>SEL_mux, O=>output_row_19);

	mux_row_20: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_20_0, I1=>output_MAC_20_1, I2=>output_MAC_20_2, I3=>output_MAC_20_3, I4=>output_MAC_20_4, I5=>output_MAC_20_5, I6=>output_MAC_20_6, I7=>output_MAC_20_7, I8=>output_MAC_20_8, I9=>output_MAC_20_9, I10=>output_MAC_20_10, I11=>output_MAC_20_11, I12=>output_MAC_20_12, I13=>output_MAC_20_13, I14=>output_MAC_20_14, I15=>output_MAC_20_15, 
		SEL_mux=>SEL_mux, O=>output_row_20);

	mux_row_21: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_21_0, I1=>output_MAC_21_1, I2=>output_MAC_21_2, I3=>output_MAC_21_3, I4=>output_MAC_21_4, I5=>output_MAC_21_5, I6=>output_MAC_21_6, I7=>output_MAC_21_7, I8=>output_MAC_21_8, I9=>output_MAC_21_9, I10=>output_MAC_21_10, I11=>output_MAC_21_11, I12=>output_MAC_21_12, I13=>output_MAC_21_13, I14=>output_MAC_21_14, I15=>output_MAC_21_15, 
		SEL_mux=>SEL_mux, O=>output_row_21);

	mux_row_22: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_22_0, I1=>output_MAC_22_1, I2=>output_MAC_22_2, I3=>output_MAC_22_3, I4=>output_MAC_22_4, I5=>output_MAC_22_5, I6=>output_MAC_22_6, I7=>output_MAC_22_7, I8=>output_MAC_22_8, I9=>output_MAC_22_9, I10=>output_MAC_22_10, I11=>output_MAC_22_11, I12=>output_MAC_22_12, I13=>output_MAC_22_13, I14=>output_MAC_22_14, I15=>output_MAC_22_15, 
		SEL_mux=>SEL_mux, O=>output_row_22);

	mux_row_23: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_23_0, I1=>output_MAC_23_1, I2=>output_MAC_23_2, I3=>output_MAC_23_3, I4=>output_MAC_23_4, I5=>output_MAC_23_5, I6=>output_MAC_23_6, I7=>output_MAC_23_7, I8=>output_MAC_23_8, I9=>output_MAC_23_9, I10=>output_MAC_23_10, I11=>output_MAC_23_11, I12=>output_MAC_23_12, I13=>output_MAC_23_13, I14=>output_MAC_23_14, I15=>output_MAC_23_15, 
		SEL_mux=>SEL_mux, O=>output_row_23);

	mux_row_24: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_24_0, I1=>output_MAC_24_1, I2=>output_MAC_24_2, I3=>output_MAC_24_3, I4=>output_MAC_24_4, I5=>output_MAC_24_5, I6=>output_MAC_24_6, I7=>output_MAC_24_7, I8=>output_MAC_24_8, I9=>output_MAC_24_9, I10=>output_MAC_24_10, I11=>output_MAC_24_11, I12=>output_MAC_24_12, I13=>output_MAC_24_13, I14=>output_MAC_24_14, I15=>output_MAC_24_15, 
		SEL_mux=>SEL_mux, O=>output_row_24);

	mux_row_25: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_25_0, I1=>output_MAC_25_1, I2=>output_MAC_25_2, I3=>output_MAC_25_3, I4=>output_MAC_25_4, I5=>output_MAC_25_5, I6=>output_MAC_25_6, I7=>output_MAC_25_7, I8=>output_MAC_25_8, I9=>output_MAC_25_9, I10=>output_MAC_25_10, I11=>output_MAC_25_11, I12=>output_MAC_25_12, I13=>output_MAC_25_13, I14=>output_MAC_25_14, I15=>output_MAC_25_15, 
		SEL_mux=>SEL_mux, O=>output_row_25);

	mux_row_26: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_26_0, I1=>output_MAC_26_1, I2=>output_MAC_26_2, I3=>output_MAC_26_3, I4=>output_MAC_26_4, I5=>output_MAC_26_5, I6=>output_MAC_26_6, I7=>output_MAC_26_7, I8=>output_MAC_26_8, I9=>output_MAC_26_9, I10=>output_MAC_26_10, I11=>output_MAC_26_11, I12=>output_MAC_26_12, I13=>output_MAC_26_13, I14=>output_MAC_26_14, I15=>output_MAC_26_15, 
		SEL_mux=>SEL_mux, O=>output_row_26);

	mux_row_27: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_27_0, I1=>output_MAC_27_1, I2=>output_MAC_27_2, I3=>output_MAC_27_3, I4=>output_MAC_27_4, I5=>output_MAC_27_5, I6=>output_MAC_27_6, I7=>output_MAC_27_7, I8=>output_MAC_27_8, I9=>output_MAC_27_9, I10=>output_MAC_27_10, I11=>output_MAC_27_11, I12=>output_MAC_27_12, I13=>output_MAC_27_13, I14=>output_MAC_27_14, I15=>output_MAC_27_15, 
		SEL_mux=>SEL_mux, O=>output_row_27);

	mux_row_28: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_28_0, I1=>output_MAC_28_1, I2=>output_MAC_28_2, I3=>output_MAC_28_3, I4=>output_MAC_28_4, I5=>output_MAC_28_5, I6=>output_MAC_28_6, I7=>output_MAC_28_7, I8=>output_MAC_28_8, I9=>output_MAC_28_9, I10=>output_MAC_28_10, I11=>output_MAC_28_11, I12=>output_MAC_28_12, I13=>output_MAC_28_13, I14=>output_MAC_28_14, I15=>output_MAC_28_15, 
		SEL_mux=>SEL_mux, O=>output_row_28);

	mux_row_29: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_29_0, I1=>output_MAC_29_1, I2=>output_MAC_29_2, I3=>output_MAC_29_3, I4=>output_MAC_29_4, I5=>output_MAC_29_5, I6=>output_MAC_29_6, I7=>output_MAC_29_7, I8=>output_MAC_29_8, I9=>output_MAC_29_9, I10=>output_MAC_29_10, I11=>output_MAC_29_11, I12=>output_MAC_29_12, I13=>output_MAC_29_13, I14=>output_MAC_29_14, I15=>output_MAC_29_15, 
		SEL_mux=>SEL_mux, O=>output_row_29);

	mux_row_30: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_30_0, I1=>output_MAC_30_1, I2=>output_MAC_30_2, I3=>output_MAC_30_3, I4=>output_MAC_30_4, I5=>output_MAC_30_5, I6=>output_MAC_30_6, I7=>output_MAC_30_7, I8=>output_MAC_30_8, I9=>output_MAC_30_9, I10=>output_MAC_30_10, I11=>output_MAC_30_11, I12=>output_MAC_30_12, I13=>output_MAC_30_13, I14=>output_MAC_30_14, I15=>output_MAC_30_15, 
		SEL_mux=>SEL_mux, O=>output_row_30);

	mux_row_31: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_31_0, I1=>output_MAC_31_1, I2=>output_MAC_31_2, I3=>output_MAC_31_3, I4=>output_MAC_31_4, I5=>output_MAC_31_5, I6=>output_MAC_31_6, I7=>output_MAC_31_7, I8=>output_MAC_31_8, I9=>output_MAC_31_9, I10=>output_MAC_31_10, I11=>output_MAC_31_11, I12=>output_MAC_31_12, I13=>output_MAC_31_13, I14=>output_MAC_31_14, I15=>output_MAC_31_15, 
		SEL_mux=>SEL_mux, O=>output_row_31);

	mux_row_32: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_32_0, I1=>output_MAC_32_1, I2=>output_MAC_32_2, I3=>output_MAC_32_3, I4=>output_MAC_32_4, I5=>output_MAC_32_5, I6=>output_MAC_32_6, I7=>output_MAC_32_7, I8=>output_MAC_32_8, I9=>output_MAC_32_9, I10=>output_MAC_32_10, I11=>output_MAC_32_11, I12=>output_MAC_32_12, I13=>output_MAC_32_13, I14=>output_MAC_32_14, I15=>output_MAC_32_15, 
		SEL_mux=>SEL_mux, O=>output_row_32);

	mux_row_33: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_33_0, I1=>output_MAC_33_1, I2=>output_MAC_33_2, I3=>output_MAC_33_3, I4=>output_MAC_33_4, I5=>output_MAC_33_5, I6=>output_MAC_33_6, I7=>output_MAC_33_7, I8=>output_MAC_33_8, I9=>output_MAC_33_9, I10=>output_MAC_33_10, I11=>output_MAC_33_11, I12=>output_MAC_33_12, I13=>output_MAC_33_13, I14=>output_MAC_33_14, I15=>output_MAC_33_15, 
		SEL_mux=>SEL_mux, O=>output_row_33);

	mux_row_34: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_34_0, I1=>output_MAC_34_1, I2=>output_MAC_34_2, I3=>output_MAC_34_3, I4=>output_MAC_34_4, I5=>output_MAC_34_5, I6=>output_MAC_34_6, I7=>output_MAC_34_7, I8=>output_MAC_34_8, I9=>output_MAC_34_9, I10=>output_MAC_34_10, I11=>output_MAC_34_11, I12=>output_MAC_34_12, I13=>output_MAC_34_13, I14=>output_MAC_34_14, I15=>output_MAC_34_15, 
		SEL_mux=>SEL_mux, O=>output_row_34);

	mux_row_35: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_35_0, I1=>output_MAC_35_1, I2=>output_MAC_35_2, I3=>output_MAC_35_3, I4=>output_MAC_35_4, I5=>output_MAC_35_5, I6=>output_MAC_35_6, I7=>output_MAC_35_7, I8=>output_MAC_35_8, I9=>output_MAC_35_9, I10=>output_MAC_35_10, I11=>output_MAC_35_11, I12=>output_MAC_35_12, I13=>output_MAC_35_13, I14=>output_MAC_35_14, I15=>output_MAC_35_15, 
		SEL_mux=>SEL_mux, O=>output_row_35);

	mux_row_36: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_36_0, I1=>output_MAC_36_1, I2=>output_MAC_36_2, I3=>output_MAC_36_3, I4=>output_MAC_36_4, I5=>output_MAC_36_5, I6=>output_MAC_36_6, I7=>output_MAC_36_7, I8=>output_MAC_36_8, I9=>output_MAC_36_9, I10=>output_MAC_36_10, I11=>output_MAC_36_11, I12=>output_MAC_36_12, I13=>output_MAC_36_13, I14=>output_MAC_36_14, I15=>output_MAC_36_15, 
		SEL_mux=>SEL_mux, O=>output_row_36);

	mux_row_37: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_37_0, I1=>output_MAC_37_1, I2=>output_MAC_37_2, I3=>output_MAC_37_3, I4=>output_MAC_37_4, I5=>output_MAC_37_5, I6=>output_MAC_37_6, I7=>output_MAC_37_7, I8=>output_MAC_37_8, I9=>output_MAC_37_9, I10=>output_MAC_37_10, I11=>output_MAC_37_11, I12=>output_MAC_37_12, I13=>output_MAC_37_13, I14=>output_MAC_37_14, I15=>output_MAC_37_15, 
		SEL_mux=>SEL_mux, O=>output_row_37);

	mux_row_38: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_38_0, I1=>output_MAC_38_1, I2=>output_MAC_38_2, I3=>output_MAC_38_3, I4=>output_MAC_38_4, I5=>output_MAC_38_5, I6=>output_MAC_38_6, I7=>output_MAC_38_7, I8=>output_MAC_38_8, I9=>output_MAC_38_9, I10=>output_MAC_38_10, I11=>output_MAC_38_11, I12=>output_MAC_38_12, I13=>output_MAC_38_13, I14=>output_MAC_38_14, I15=>output_MAC_38_15, 
		SEL_mux=>SEL_mux, O=>output_row_38);

	mux_row_39: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_39_0, I1=>output_MAC_39_1, I2=>output_MAC_39_2, I3=>output_MAC_39_3, I4=>output_MAC_39_4, I5=>output_MAC_39_5, I6=>output_MAC_39_6, I7=>output_MAC_39_7, I8=>output_MAC_39_8, I9=>output_MAC_39_9, I10=>output_MAC_39_10, I11=>output_MAC_39_11, I12=>output_MAC_39_12, I13=>output_MAC_39_13, I14=>output_MAC_39_14, I15=>output_MAC_39_15, 
		SEL_mux=>SEL_mux, O=>output_row_39);

	mux_row_40: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_40_0, I1=>output_MAC_40_1, I2=>output_MAC_40_2, I3=>output_MAC_40_3, I4=>output_MAC_40_4, I5=>output_MAC_40_5, I6=>output_MAC_40_6, I7=>output_MAC_40_7, I8=>output_MAC_40_8, I9=>output_MAC_40_9, I10=>output_MAC_40_10, I11=>output_MAC_40_11, I12=>output_MAC_40_12, I13=>output_MAC_40_13, I14=>output_MAC_40_14, I15=>output_MAC_40_15, 
		SEL_mux=>SEL_mux, O=>output_row_40);

	mux_row_41: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_41_0, I1=>output_MAC_41_1, I2=>output_MAC_41_2, I3=>output_MAC_41_3, I4=>output_MAC_41_4, I5=>output_MAC_41_5, I6=>output_MAC_41_6, I7=>output_MAC_41_7, I8=>output_MAC_41_8, I9=>output_MAC_41_9, I10=>output_MAC_41_10, I11=>output_MAC_41_11, I12=>output_MAC_41_12, I13=>output_MAC_41_13, I14=>output_MAC_41_14, I15=>output_MAC_41_15, 
		SEL_mux=>SEL_mux, O=>output_row_41);

	mux_row_42: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_42_0, I1=>output_MAC_42_1, I2=>output_MAC_42_2, I3=>output_MAC_42_3, I4=>output_MAC_42_4, I5=>output_MAC_42_5, I6=>output_MAC_42_6, I7=>output_MAC_42_7, I8=>output_MAC_42_8, I9=>output_MAC_42_9, I10=>output_MAC_42_10, I11=>output_MAC_42_11, I12=>output_MAC_42_12, I13=>output_MAC_42_13, I14=>output_MAC_42_14, I15=>output_MAC_42_15, 
		SEL_mux=>SEL_mux, O=>output_row_42);

	mux_row_43: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_43_0, I1=>output_MAC_43_1, I2=>output_MAC_43_2, I3=>output_MAC_43_3, I4=>output_MAC_43_4, I5=>output_MAC_43_5, I6=>output_MAC_43_6, I7=>output_MAC_43_7, I8=>output_MAC_43_8, I9=>output_MAC_43_9, I10=>output_MAC_43_10, I11=>output_MAC_43_11, I12=>output_MAC_43_12, I13=>output_MAC_43_13, I14=>output_MAC_43_14, I15=>output_MAC_43_15, 
		SEL_mux=>SEL_mux, O=>output_row_43);

	mux_row_44: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_44_0, I1=>output_MAC_44_1, I2=>output_MAC_44_2, I3=>output_MAC_44_3, I4=>output_MAC_44_4, I5=>output_MAC_44_5, I6=>output_MAC_44_6, I7=>output_MAC_44_7, I8=>output_MAC_44_8, I9=>output_MAC_44_9, I10=>output_MAC_44_10, I11=>output_MAC_44_11, I12=>output_MAC_44_12, I13=>output_MAC_44_13, I14=>output_MAC_44_14, I15=>output_MAC_44_15, 
		SEL_mux=>SEL_mux, O=>output_row_44);

	mux_row_45: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_45_0, I1=>output_MAC_45_1, I2=>output_MAC_45_2, I3=>output_MAC_45_3, I4=>output_MAC_45_4, I5=>output_MAC_45_5, I6=>output_MAC_45_6, I7=>output_MAC_45_7, I8=>output_MAC_45_8, I9=>output_MAC_45_9, I10=>output_MAC_45_10, I11=>output_MAC_45_11, I12=>output_MAC_45_12, I13=>output_MAC_45_13, I14=>output_MAC_45_14, I15=>output_MAC_45_15, 
		SEL_mux=>SEL_mux, O=>output_row_45);

	mux_row_46: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_46_0, I1=>output_MAC_46_1, I2=>output_MAC_46_2, I3=>output_MAC_46_3, I4=>output_MAC_46_4, I5=>output_MAC_46_5, I6=>output_MAC_46_6, I7=>output_MAC_46_7, I8=>output_MAC_46_8, I9=>output_MAC_46_9, I10=>output_MAC_46_10, I11=>output_MAC_46_11, I12=>output_MAC_46_12, I13=>output_MAC_46_13, I14=>output_MAC_46_14, I15=>output_MAC_46_15, 
		SEL_mux=>SEL_mux, O=>output_row_46);

	mux_row_47: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_47_0, I1=>output_MAC_47_1, I2=>output_MAC_47_2, I3=>output_MAC_47_3, I4=>output_MAC_47_4, I5=>output_MAC_47_5, I6=>output_MAC_47_6, I7=>output_MAC_47_7, I8=>output_MAC_47_8, I9=>output_MAC_47_9, I10=>output_MAC_47_10, I11=>output_MAC_47_11, I12=>output_MAC_47_12, I13=>output_MAC_47_13, I14=>output_MAC_47_14, I15=>output_MAC_47_15, 
		SEL_mux=>SEL_mux, O=>output_row_47);

	mux_row_48: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_48_0, I1=>output_MAC_48_1, I2=>output_MAC_48_2, I3=>output_MAC_48_3, I4=>output_MAC_48_4, I5=>output_MAC_48_5, I6=>output_MAC_48_6, I7=>output_MAC_48_7, I8=>output_MAC_48_8, I9=>output_MAC_48_9, I10=>output_MAC_48_10, I11=>output_MAC_48_11, I12=>output_MAC_48_12, I13=>output_MAC_48_13, I14=>output_MAC_48_14, I15=>output_MAC_48_15, 
		SEL_mux=>SEL_mux, O=>output_row_48);

	mux_row_49: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_49_0, I1=>output_MAC_49_1, I2=>output_MAC_49_2, I3=>output_MAC_49_3, I4=>output_MAC_49_4, I5=>output_MAC_49_5, I6=>output_MAC_49_6, I7=>output_MAC_49_7, I8=>output_MAC_49_8, I9=>output_MAC_49_9, I10=>output_MAC_49_10, I11=>output_MAC_49_11, I12=>output_MAC_49_12, I13=>output_MAC_49_13, I14=>output_MAC_49_14, I15=>output_MAC_49_15, 
		SEL_mux=>SEL_mux, O=>output_row_49);

	mux_row_50: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_50_0, I1=>output_MAC_50_1, I2=>output_MAC_50_2, I3=>output_MAC_50_3, I4=>output_MAC_50_4, I5=>output_MAC_50_5, I6=>output_MAC_50_6, I7=>output_MAC_50_7, I8=>output_MAC_50_8, I9=>output_MAC_50_9, I10=>output_MAC_50_10, I11=>output_MAC_50_11, I12=>output_MAC_50_12, I13=>output_MAC_50_13, I14=>output_MAC_50_14, I15=>output_MAC_50_15, 
		SEL_mux=>SEL_mux, O=>output_row_50);

	mux_row_51: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_51_0, I1=>output_MAC_51_1, I2=>output_MAC_51_2, I3=>output_MAC_51_3, I4=>output_MAC_51_4, I5=>output_MAC_51_5, I6=>output_MAC_51_6, I7=>output_MAC_51_7, I8=>output_MAC_51_8, I9=>output_MAC_51_9, I10=>output_MAC_51_10, I11=>output_MAC_51_11, I12=>output_MAC_51_12, I13=>output_MAC_51_13, I14=>output_MAC_51_14, I15=>output_MAC_51_15, 
		SEL_mux=>SEL_mux, O=>output_row_51);

	mux_row_52: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_52_0, I1=>output_MAC_52_1, I2=>output_MAC_52_2, I3=>output_MAC_52_3, I4=>output_MAC_52_4, I5=>output_MAC_52_5, I6=>output_MAC_52_6, I7=>output_MAC_52_7, I8=>output_MAC_52_8, I9=>output_MAC_52_9, I10=>output_MAC_52_10, I11=>output_MAC_52_11, I12=>output_MAC_52_12, I13=>output_MAC_52_13, I14=>output_MAC_52_14, I15=>output_MAC_52_15, 
		SEL_mux=>SEL_mux, O=>output_row_52);

	mux_row_53: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_53_0, I1=>output_MAC_53_1, I2=>output_MAC_53_2, I3=>output_MAC_53_3, I4=>output_MAC_53_4, I5=>output_MAC_53_5, I6=>output_MAC_53_6, I7=>output_MAC_53_7, I8=>output_MAC_53_8, I9=>output_MAC_53_9, I10=>output_MAC_53_10, I11=>output_MAC_53_11, I12=>output_MAC_53_12, I13=>output_MAC_53_13, I14=>output_MAC_53_14, I15=>output_MAC_53_15, 
		SEL_mux=>SEL_mux, O=>output_row_53);

	mux_row_54: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_54_0, I1=>output_MAC_54_1, I2=>output_MAC_54_2, I3=>output_MAC_54_3, I4=>output_MAC_54_4, I5=>output_MAC_54_5, I6=>output_MAC_54_6, I7=>output_MAC_54_7, I8=>output_MAC_54_8, I9=>output_MAC_54_9, I10=>output_MAC_54_10, I11=>output_MAC_54_11, I12=>output_MAC_54_12, I13=>output_MAC_54_13, I14=>output_MAC_54_14, I15=>output_MAC_54_15, 
		SEL_mux=>SEL_mux, O=>output_row_54);

	mux_row_55: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_55_0, I1=>output_MAC_55_1, I2=>output_MAC_55_2, I3=>output_MAC_55_3, I4=>output_MAC_55_4, I5=>output_MAC_55_5, I6=>output_MAC_55_6, I7=>output_MAC_55_7, I8=>output_MAC_55_8, I9=>output_MAC_55_9, I10=>output_MAC_55_10, I11=>output_MAC_55_11, I12=>output_MAC_55_12, I13=>output_MAC_55_13, I14=>output_MAC_55_14, I15=>output_MAC_55_15, 
		SEL_mux=>SEL_mux, O=>output_row_55);

	mux_row_56: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_56_0, I1=>output_MAC_56_1, I2=>output_MAC_56_2, I3=>output_MAC_56_3, I4=>output_MAC_56_4, I5=>output_MAC_56_5, I6=>output_MAC_56_6, I7=>output_MAC_56_7, I8=>output_MAC_56_8, I9=>output_MAC_56_9, I10=>output_MAC_56_10, I11=>output_MAC_56_11, I12=>output_MAC_56_12, I13=>output_MAC_56_13, I14=>output_MAC_56_14, I15=>output_MAC_56_15, 
		SEL_mux=>SEL_mux, O=>output_row_56);

	mux_row_57: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_57_0, I1=>output_MAC_57_1, I2=>output_MAC_57_2, I3=>output_MAC_57_3, I4=>output_MAC_57_4, I5=>output_MAC_57_5, I6=>output_MAC_57_6, I7=>output_MAC_57_7, I8=>output_MAC_57_8, I9=>output_MAC_57_9, I10=>output_MAC_57_10, I11=>output_MAC_57_11, I12=>output_MAC_57_12, I13=>output_MAC_57_13, I14=>output_MAC_57_14, I15=>output_MAC_57_15, 
		SEL_mux=>SEL_mux, O=>output_row_57);

	mux_row_58: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_58_0, I1=>output_MAC_58_1, I2=>output_MAC_58_2, I3=>output_MAC_58_3, I4=>output_MAC_58_4, I5=>output_MAC_58_5, I6=>output_MAC_58_6, I7=>output_MAC_58_7, I8=>output_MAC_58_8, I9=>output_MAC_58_9, I10=>output_MAC_58_10, I11=>output_MAC_58_11, I12=>output_MAC_58_12, I13=>output_MAC_58_13, I14=>output_MAC_58_14, I15=>output_MAC_58_15, 
		SEL_mux=>SEL_mux, O=>output_row_58);

	mux_row_59: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_59_0, I1=>output_MAC_59_1, I2=>output_MAC_59_2, I3=>output_MAC_59_3, I4=>output_MAC_59_4, I5=>output_MAC_59_5, I6=>output_MAC_59_6, I7=>output_MAC_59_7, I8=>output_MAC_59_8, I9=>output_MAC_59_9, I10=>output_MAC_59_10, I11=>output_MAC_59_11, I12=>output_MAC_59_12, I13=>output_MAC_59_13, I14=>output_MAC_59_14, I15=>output_MAC_59_15, 
		SEL_mux=>SEL_mux, O=>output_row_59);

	mux_row_60: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_60_0, I1=>output_MAC_60_1, I2=>output_MAC_60_2, I3=>output_MAC_60_3, I4=>output_MAC_60_4, I5=>output_MAC_60_5, I6=>output_MAC_60_6, I7=>output_MAC_60_7, I8=>output_MAC_60_8, I9=>output_MAC_60_9, I10=>output_MAC_60_10, I11=>output_MAC_60_11, I12=>output_MAC_60_12, I13=>output_MAC_60_13, I14=>output_MAC_60_14, I15=>output_MAC_60_15, 
		SEL_mux=>SEL_mux, O=>output_row_60);

	mux_row_61: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_61_0, I1=>output_MAC_61_1, I2=>output_MAC_61_2, I3=>output_MAC_61_3, I4=>output_MAC_61_4, I5=>output_MAC_61_5, I6=>output_MAC_61_6, I7=>output_MAC_61_7, I8=>output_MAC_61_8, I9=>output_MAC_61_9, I10=>output_MAC_61_10, I11=>output_MAC_61_11, I12=>output_MAC_61_12, I13=>output_MAC_61_13, I14=>output_MAC_61_14, I15=>output_MAC_61_15, 
		SEL_mux=>SEL_mux, O=>output_row_61);

	mux_row_62: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_62_0, I1=>output_MAC_62_1, I2=>output_MAC_62_2, I3=>output_MAC_62_3, I4=>output_MAC_62_4, I5=>output_MAC_62_5, I6=>output_MAC_62_6, I7=>output_MAC_62_7, I8=>output_MAC_62_8, I9=>output_MAC_62_9, I10=>output_MAC_62_10, I11=>output_MAC_62_11, I12=>output_MAC_62_12, I13=>output_MAC_62_13, I14=>output_MAC_62_14, I15=>output_MAC_62_15, 
		SEL_mux=>SEL_mux, O=>output_row_62);

	mux_row_63: mux_16to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_63_0, I1=>output_MAC_63_1, I2=>output_MAC_63_2, I3=>output_MAC_63_3, I4=>output_MAC_63_4, I5=>output_MAC_63_5, I6=>output_MAC_63_6, I7=>output_MAC_63_7, I8=>output_MAC_63_8, I9=>output_MAC_63_9, I10=>output_MAC_63_10, I11=>output_MAC_63_11, I12=>output_MAC_63_12, I13=>output_MAC_63_13, I14=>output_MAC_63_14, I15=>output_MAC_63_15, 
		SEL_mux=>SEL_mux, O=>output_row_63);


END behaviour;
