
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MAC_128x32_8_reg IS
PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7, input_row_8, input_row_9, 
	input_row_10, input_row_11, input_row_12, input_row_13, input_row_14, input_row_15, input_row_16, input_row_17, input_row_18, input_row_19, 
	input_row_20, input_row_21, input_row_22, input_row_23, input_row_24, input_row_25, input_row_26, input_row_27, input_row_28, input_row_29, 
	input_row_30, input_row_31, input_row_32, input_row_33, input_row_34, input_row_35, input_row_36, input_row_37, input_row_38, input_row_39, 
	input_row_40, input_row_41, input_row_42, input_row_43, input_row_44, input_row_45, input_row_46, input_row_47, input_row_48, input_row_49, 
	input_row_50, input_row_51, input_row_52, input_row_53, input_row_54, input_row_55, input_row_56, input_row_57, input_row_58, input_row_59, 
	input_row_60, input_row_61, input_row_62, input_row_63, input_row_64, input_row_65, input_row_66, input_row_67, input_row_68, input_row_69, 
	input_row_70, input_row_71, input_row_72, input_row_73, input_row_74, input_row_75, input_row_76, input_row_77, input_row_78, input_row_79, 
	input_row_80, input_row_81, input_row_82, input_row_83, input_row_84, input_row_85, input_row_86, input_row_87, input_row_88, input_row_89, 
	input_row_90, input_row_91, input_row_92, input_row_93, input_row_94, input_row_95, input_row_96, input_row_97, input_row_98, input_row_99, 
	input_row_100, input_row_101, input_row_102, input_row_103, input_row_104, input_row_105, input_row_106, input_row_107, input_row_108, input_row_109, 
	input_row_110, input_row_111, input_row_112, input_row_113, input_row_114, input_row_115, input_row_116, input_row_117, input_row_118, input_row_119, 
	input_row_120, input_row_121, input_row_122, input_row_123, input_row_124, input_row_125, input_row_126, input_row_127: IN STD_LOGIC_VECTOR(7 downto 0);
	input_col_0, input_col_1, input_col_2, input_col_3, input_col_4, input_col_5, input_col_6, input_col_7, input_col_8, input_col_9, 
	input_col_10, input_col_11, input_col_12, input_col_13, input_col_14, input_col_15, input_col_16, input_col_17, input_col_18, input_col_19, 
	input_col_20, input_col_21, input_col_22, input_col_23, input_col_24, input_col_25, input_col_26, input_col_27, input_col_28, input_col_29, 
	input_col_30, input_col_31: IN STD_LOGIC_VECTOR(7 downto 0);
	SEL_mux: IN STD_LOGIC_VECTOR(4 downto 0);
	CLK, RST_n, ENABLE : IN STD_LOGIC;
	output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7, output_row_8, output_row_9, 
	output_row_10, output_row_11, output_row_12, output_row_13, output_row_14, output_row_15, output_row_16, output_row_17, output_row_18, output_row_19, 
	output_row_20, output_row_21, output_row_22, output_row_23, output_row_24, output_row_25, output_row_26, output_row_27, output_row_28, output_row_29, 
	output_row_30, output_row_31, output_row_32, output_row_33, output_row_34, output_row_35, output_row_36, output_row_37, output_row_38, output_row_39, 
	output_row_40, output_row_41, output_row_42, output_row_43, output_row_44, output_row_45, output_row_46, output_row_47, output_row_48, output_row_49, 
	output_row_50, output_row_51, output_row_52, output_row_53, output_row_54, output_row_55, output_row_56, output_row_57, output_row_58, output_row_59, 
	output_row_60, output_row_61, output_row_62, output_row_63, output_row_64, output_row_65, output_row_66, output_row_67, output_row_68, output_row_69, 
	output_row_70, output_row_71, output_row_72, output_row_73, output_row_74, output_row_75, output_row_76, output_row_77, output_row_78, output_row_79, 
	output_row_80, output_row_81, output_row_82, output_row_83, output_row_84, output_row_85, output_row_86, output_row_87, output_row_88, output_row_89, 
	output_row_90, output_row_91, output_row_92, output_row_93, output_row_94, output_row_95, output_row_96, output_row_97, output_row_98, output_row_99, 
	output_row_100, output_row_101, output_row_102, output_row_103, output_row_104, output_row_105, output_row_106, output_row_107, output_row_108, output_row_109, 
	output_row_110, output_row_111, output_row_112, output_row_113, output_row_114, output_row_115, output_row_116, output_row_117, output_row_118, output_row_119, 
	output_row_120, output_row_121, output_row_122, output_row_123, output_row_124, output_row_125, output_row_126, output_row_127: OUT STD_LOGIC_VECTOR(31 downto 0)
);
END MAC_128x32_8_reg;

ARCHITECTURE behaviour OF  MAC_128x32_8_reg IS

	COMPONENT MAC IS
	GENERIC (data_size : POSITIVE := 2; 
	acc_size: POSITIVE := 16	);
	PORT( data_in_A, data_in_B  : IN STD_LOGIC_VECTOR(data_size-1 downto 0);
		CLK, RST_n, ENABLE 	: IN STD_LOGIC;
		data_out    			: OUT STD_LOGIC_VECTOR(acc_size-1 downto 0));
	END COMPONENT;

	COMPONENT mux_32to1_nbit IS
	GENERIC ( N : POSITIVE :=2);
	PORT(
		I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, 
		I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, 
		I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, 
		I30, I31: IN STD_LOGIC_VECTOR(N-1 downto 0);
		SEL_mux  : IN STD_LOGIC_VECTOR(4 downto 0);
		O    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
	END COMPONENT;

	COMPONENT regnbit IS
	GENERIC ( N : POSITIVE := 2);
	PORT(
		D    : IN STD_LOGIC_VECTOR(N-1 downto 0);
		CLK, RST_n, ENABLE : IN STD_LOGIC;
		Q    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
	END COMPONENT;

	COMPONENT ff IS
	PORT(
		D    : IN STD_LOGIC;
		CLK, RST_n, ENABLE : IN STD_LOGIC;
		Q    : OUT STD_LOGIC
	);
	END COMPONENT;

	SIGNAL reg_input_row_0, reg_input_row_1, reg_input_row_2, reg_input_row_3, reg_input_row_4, reg_input_row_5, reg_input_row_6, reg_input_row_7, reg_input_row_8, reg_input_row_9, 
		reg_input_row_10, reg_input_row_11, reg_input_row_12, reg_input_row_13, reg_input_row_14, reg_input_row_15, reg_input_row_16, reg_input_row_17, reg_input_row_18, reg_input_row_19, 
		reg_input_row_20, reg_input_row_21, reg_input_row_22, reg_input_row_23, reg_input_row_24, reg_input_row_25, reg_input_row_26, reg_input_row_27, reg_input_row_28, reg_input_row_29, 
		reg_input_row_30, reg_input_row_31, reg_input_row_32, reg_input_row_33, reg_input_row_34, reg_input_row_35, reg_input_row_36, reg_input_row_37, reg_input_row_38, reg_input_row_39, 
		reg_input_row_40, reg_input_row_41, reg_input_row_42, reg_input_row_43, reg_input_row_44, reg_input_row_45, reg_input_row_46, reg_input_row_47, reg_input_row_48, reg_input_row_49, 
		reg_input_row_50, reg_input_row_51, reg_input_row_52, reg_input_row_53, reg_input_row_54, reg_input_row_55, reg_input_row_56, reg_input_row_57, reg_input_row_58, reg_input_row_59, 
		reg_input_row_60, reg_input_row_61, reg_input_row_62, reg_input_row_63, reg_input_row_64, reg_input_row_65, reg_input_row_66, reg_input_row_67, reg_input_row_68, reg_input_row_69, 
		reg_input_row_70, reg_input_row_71, reg_input_row_72, reg_input_row_73, reg_input_row_74, reg_input_row_75, reg_input_row_76, reg_input_row_77, reg_input_row_78, reg_input_row_79, 
		reg_input_row_80, reg_input_row_81, reg_input_row_82, reg_input_row_83, reg_input_row_84, reg_input_row_85, reg_input_row_86, reg_input_row_87, reg_input_row_88, reg_input_row_89, 
		reg_input_row_90, reg_input_row_91, reg_input_row_92, reg_input_row_93, reg_input_row_94, reg_input_row_95, reg_input_row_96, reg_input_row_97, reg_input_row_98, reg_input_row_99, 
		reg_input_row_100, reg_input_row_101, reg_input_row_102, reg_input_row_103, reg_input_row_104, reg_input_row_105, reg_input_row_106, reg_input_row_107, reg_input_row_108, reg_input_row_109, 
		reg_input_row_110, reg_input_row_111, reg_input_row_112, reg_input_row_113, reg_input_row_114, reg_input_row_115, reg_input_row_116, reg_input_row_117, reg_input_row_118, reg_input_row_119, 
		reg_input_row_120, reg_input_row_121, reg_input_row_122, reg_input_row_123, reg_input_row_124, reg_input_row_125, reg_input_row_126, reg_input_row_127: STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL reg_input_col_0, reg_input_col_1, reg_input_col_2, reg_input_col_3, reg_input_col_4, reg_input_col_5, reg_input_col_6, reg_input_col_7, reg_input_col_8, reg_input_col_9, 
		reg_input_col_10, reg_input_col_11, reg_input_col_12, reg_input_col_13, reg_input_col_14, reg_input_col_15, reg_input_col_16, reg_input_col_17, reg_input_col_18, reg_input_col_19, 
		reg_input_col_20, reg_input_col_21, reg_input_col_22, reg_input_col_23, reg_input_col_24, reg_input_col_25, reg_input_col_26, reg_input_col_27, reg_input_col_28, reg_input_col_29, 
		reg_input_col_30, reg_input_col_31: STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL reg_SEL_mux: STD_LOGIC_VECTOR(4 downto 0);
	SIGNAL reg_ENABLE_in, reg_ENABLE_out : STD_LOGIC;
	SIGNAL reg_output_row_0, reg_output_row_1, reg_output_row_2, reg_output_row_3, reg_output_row_4, reg_output_row_5, reg_output_row_6, reg_output_row_7, reg_output_row_8, reg_output_row_9, 
		reg_output_row_10, reg_output_row_11, reg_output_row_12, reg_output_row_13, reg_output_row_14, reg_output_row_15, reg_output_row_16, reg_output_row_17, reg_output_row_18, reg_output_row_19, 
		reg_output_row_20, reg_output_row_21, reg_output_row_22, reg_output_row_23, reg_output_row_24, reg_output_row_25, reg_output_row_26, reg_output_row_27, reg_output_row_28, reg_output_row_29, 
		reg_output_row_30, reg_output_row_31, reg_output_row_32, reg_output_row_33, reg_output_row_34, reg_output_row_35, reg_output_row_36, reg_output_row_37, reg_output_row_38, reg_output_row_39, 
		reg_output_row_40, reg_output_row_41, reg_output_row_42, reg_output_row_43, reg_output_row_44, reg_output_row_45, reg_output_row_46, reg_output_row_47, reg_output_row_48, reg_output_row_49, 
		reg_output_row_50, reg_output_row_51, reg_output_row_52, reg_output_row_53, reg_output_row_54, reg_output_row_55, reg_output_row_56, reg_output_row_57, reg_output_row_58, reg_output_row_59, 
		reg_output_row_60, reg_output_row_61, reg_output_row_62, reg_output_row_63, reg_output_row_64, reg_output_row_65, reg_output_row_66, reg_output_row_67, reg_output_row_68, reg_output_row_69, 
		reg_output_row_70, reg_output_row_71, reg_output_row_72, reg_output_row_73, reg_output_row_74, reg_output_row_75, reg_output_row_76, reg_output_row_77, reg_output_row_78, reg_output_row_79, 
		reg_output_row_80, reg_output_row_81, reg_output_row_82, reg_output_row_83, reg_output_row_84, reg_output_row_85, reg_output_row_86, reg_output_row_87, reg_output_row_88, reg_output_row_89, 
		reg_output_row_90, reg_output_row_91, reg_output_row_92, reg_output_row_93, reg_output_row_94, reg_output_row_95, reg_output_row_96, reg_output_row_97, reg_output_row_98, reg_output_row_99, 
		reg_output_row_100, reg_output_row_101, reg_output_row_102, reg_output_row_103, reg_output_row_104, reg_output_row_105, reg_output_row_106, reg_output_row_107, reg_output_row_108, reg_output_row_109, 
		reg_output_row_110, reg_output_row_111, reg_output_row_112, reg_output_row_113, reg_output_row_114, reg_output_row_115, reg_output_row_116, reg_output_row_117, reg_output_row_118, reg_output_row_119, 
		reg_output_row_120, reg_output_row_121, reg_output_row_122, reg_output_row_123, reg_output_row_124, reg_output_row_125, reg_output_row_126, reg_output_row_127: STD_LOGIC_VECTOR(31 downto 0);

	SIGNAL output_MAC_0_0, output_MAC_0_1, output_MAC_0_2, output_MAC_0_3, output_MAC_0_4, output_MAC_0_5, output_MAC_0_6, output_MAC_0_7, output_MAC_0_8, output_MAC_0_9, 
		output_MAC_0_10, output_MAC_0_11, output_MAC_0_12, output_MAC_0_13, output_MAC_0_14, output_MAC_0_15, output_MAC_0_16, output_MAC_0_17, output_MAC_0_18, output_MAC_0_19, 
		output_MAC_0_20, output_MAC_0_21, output_MAC_0_22, output_MAC_0_23, output_MAC_0_24, output_MAC_0_25, output_MAC_0_26, output_MAC_0_27, output_MAC_0_28, output_MAC_0_29, 
		output_MAC_0_30, output_MAC_0_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_1_0, output_MAC_1_1, output_MAC_1_2, output_MAC_1_3, output_MAC_1_4, output_MAC_1_5, output_MAC_1_6, output_MAC_1_7, output_MAC_1_8, output_MAC_1_9, 
		output_MAC_1_10, output_MAC_1_11, output_MAC_1_12, output_MAC_1_13, output_MAC_1_14, output_MAC_1_15, output_MAC_1_16, output_MAC_1_17, output_MAC_1_18, output_MAC_1_19, 
		output_MAC_1_20, output_MAC_1_21, output_MAC_1_22, output_MAC_1_23, output_MAC_1_24, output_MAC_1_25, output_MAC_1_26, output_MAC_1_27, output_MAC_1_28, output_MAC_1_29, 
		output_MAC_1_30, output_MAC_1_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_2_0, output_MAC_2_1, output_MAC_2_2, output_MAC_2_3, output_MAC_2_4, output_MAC_2_5, output_MAC_2_6, output_MAC_2_7, output_MAC_2_8, output_MAC_2_9, 
		output_MAC_2_10, output_MAC_2_11, output_MAC_2_12, output_MAC_2_13, output_MAC_2_14, output_MAC_2_15, output_MAC_2_16, output_MAC_2_17, output_MAC_2_18, output_MAC_2_19, 
		output_MAC_2_20, output_MAC_2_21, output_MAC_2_22, output_MAC_2_23, output_MAC_2_24, output_MAC_2_25, output_MAC_2_26, output_MAC_2_27, output_MAC_2_28, output_MAC_2_29, 
		output_MAC_2_30, output_MAC_2_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_3_0, output_MAC_3_1, output_MAC_3_2, output_MAC_3_3, output_MAC_3_4, output_MAC_3_5, output_MAC_3_6, output_MAC_3_7, output_MAC_3_8, output_MAC_3_9, 
		output_MAC_3_10, output_MAC_3_11, output_MAC_3_12, output_MAC_3_13, output_MAC_3_14, output_MAC_3_15, output_MAC_3_16, output_MAC_3_17, output_MAC_3_18, output_MAC_3_19, 
		output_MAC_3_20, output_MAC_3_21, output_MAC_3_22, output_MAC_3_23, output_MAC_3_24, output_MAC_3_25, output_MAC_3_26, output_MAC_3_27, output_MAC_3_28, output_MAC_3_29, 
		output_MAC_3_30, output_MAC_3_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_4_0, output_MAC_4_1, output_MAC_4_2, output_MAC_4_3, output_MAC_4_4, output_MAC_4_5, output_MAC_4_6, output_MAC_4_7, output_MAC_4_8, output_MAC_4_9, 
		output_MAC_4_10, output_MAC_4_11, output_MAC_4_12, output_MAC_4_13, output_MAC_4_14, output_MAC_4_15, output_MAC_4_16, output_MAC_4_17, output_MAC_4_18, output_MAC_4_19, 
		output_MAC_4_20, output_MAC_4_21, output_MAC_4_22, output_MAC_4_23, output_MAC_4_24, output_MAC_4_25, output_MAC_4_26, output_MAC_4_27, output_MAC_4_28, output_MAC_4_29, 
		output_MAC_4_30, output_MAC_4_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_5_0, output_MAC_5_1, output_MAC_5_2, output_MAC_5_3, output_MAC_5_4, output_MAC_5_5, output_MAC_5_6, output_MAC_5_7, output_MAC_5_8, output_MAC_5_9, 
		output_MAC_5_10, output_MAC_5_11, output_MAC_5_12, output_MAC_5_13, output_MAC_5_14, output_MAC_5_15, output_MAC_5_16, output_MAC_5_17, output_MAC_5_18, output_MAC_5_19, 
		output_MAC_5_20, output_MAC_5_21, output_MAC_5_22, output_MAC_5_23, output_MAC_5_24, output_MAC_5_25, output_MAC_5_26, output_MAC_5_27, output_MAC_5_28, output_MAC_5_29, 
		output_MAC_5_30, output_MAC_5_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_6_0, output_MAC_6_1, output_MAC_6_2, output_MAC_6_3, output_MAC_6_4, output_MAC_6_5, output_MAC_6_6, output_MAC_6_7, output_MAC_6_8, output_MAC_6_9, 
		output_MAC_6_10, output_MAC_6_11, output_MAC_6_12, output_MAC_6_13, output_MAC_6_14, output_MAC_6_15, output_MAC_6_16, output_MAC_6_17, output_MAC_6_18, output_MAC_6_19, 
		output_MAC_6_20, output_MAC_6_21, output_MAC_6_22, output_MAC_6_23, output_MAC_6_24, output_MAC_6_25, output_MAC_6_26, output_MAC_6_27, output_MAC_6_28, output_MAC_6_29, 
		output_MAC_6_30, output_MAC_6_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_7_0, output_MAC_7_1, output_MAC_7_2, output_MAC_7_3, output_MAC_7_4, output_MAC_7_5, output_MAC_7_6, output_MAC_7_7, output_MAC_7_8, output_MAC_7_9, 
		output_MAC_7_10, output_MAC_7_11, output_MAC_7_12, output_MAC_7_13, output_MAC_7_14, output_MAC_7_15, output_MAC_7_16, output_MAC_7_17, output_MAC_7_18, output_MAC_7_19, 
		output_MAC_7_20, output_MAC_7_21, output_MAC_7_22, output_MAC_7_23, output_MAC_7_24, output_MAC_7_25, output_MAC_7_26, output_MAC_7_27, output_MAC_7_28, output_MAC_7_29, 
		output_MAC_7_30, output_MAC_7_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_8_0, output_MAC_8_1, output_MAC_8_2, output_MAC_8_3, output_MAC_8_4, output_MAC_8_5, output_MAC_8_6, output_MAC_8_7, output_MAC_8_8, output_MAC_8_9, 
		output_MAC_8_10, output_MAC_8_11, output_MAC_8_12, output_MAC_8_13, output_MAC_8_14, output_MAC_8_15, output_MAC_8_16, output_MAC_8_17, output_MAC_8_18, output_MAC_8_19, 
		output_MAC_8_20, output_MAC_8_21, output_MAC_8_22, output_MAC_8_23, output_MAC_8_24, output_MAC_8_25, output_MAC_8_26, output_MAC_8_27, output_MAC_8_28, output_MAC_8_29, 
		output_MAC_8_30, output_MAC_8_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_9_0, output_MAC_9_1, output_MAC_9_2, output_MAC_9_3, output_MAC_9_4, output_MAC_9_5, output_MAC_9_6, output_MAC_9_7, output_MAC_9_8, output_MAC_9_9, 
		output_MAC_9_10, output_MAC_9_11, output_MAC_9_12, output_MAC_9_13, output_MAC_9_14, output_MAC_9_15, output_MAC_9_16, output_MAC_9_17, output_MAC_9_18, output_MAC_9_19, 
		output_MAC_9_20, output_MAC_9_21, output_MAC_9_22, output_MAC_9_23, output_MAC_9_24, output_MAC_9_25, output_MAC_9_26, output_MAC_9_27, output_MAC_9_28, output_MAC_9_29, 
		output_MAC_9_30, output_MAC_9_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_10_0, output_MAC_10_1, output_MAC_10_2, output_MAC_10_3, output_MAC_10_4, output_MAC_10_5, output_MAC_10_6, output_MAC_10_7, output_MAC_10_8, output_MAC_10_9, 
		output_MAC_10_10, output_MAC_10_11, output_MAC_10_12, output_MAC_10_13, output_MAC_10_14, output_MAC_10_15, output_MAC_10_16, output_MAC_10_17, output_MAC_10_18, output_MAC_10_19, 
		output_MAC_10_20, output_MAC_10_21, output_MAC_10_22, output_MAC_10_23, output_MAC_10_24, output_MAC_10_25, output_MAC_10_26, output_MAC_10_27, output_MAC_10_28, output_MAC_10_29, 
		output_MAC_10_30, output_MAC_10_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_11_0, output_MAC_11_1, output_MAC_11_2, output_MAC_11_3, output_MAC_11_4, output_MAC_11_5, output_MAC_11_6, output_MAC_11_7, output_MAC_11_8, output_MAC_11_9, 
		output_MAC_11_10, output_MAC_11_11, output_MAC_11_12, output_MAC_11_13, output_MAC_11_14, output_MAC_11_15, output_MAC_11_16, output_MAC_11_17, output_MAC_11_18, output_MAC_11_19, 
		output_MAC_11_20, output_MAC_11_21, output_MAC_11_22, output_MAC_11_23, output_MAC_11_24, output_MAC_11_25, output_MAC_11_26, output_MAC_11_27, output_MAC_11_28, output_MAC_11_29, 
		output_MAC_11_30, output_MAC_11_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_12_0, output_MAC_12_1, output_MAC_12_2, output_MAC_12_3, output_MAC_12_4, output_MAC_12_5, output_MAC_12_6, output_MAC_12_7, output_MAC_12_8, output_MAC_12_9, 
		output_MAC_12_10, output_MAC_12_11, output_MAC_12_12, output_MAC_12_13, output_MAC_12_14, output_MAC_12_15, output_MAC_12_16, output_MAC_12_17, output_MAC_12_18, output_MAC_12_19, 
		output_MAC_12_20, output_MAC_12_21, output_MAC_12_22, output_MAC_12_23, output_MAC_12_24, output_MAC_12_25, output_MAC_12_26, output_MAC_12_27, output_MAC_12_28, output_MAC_12_29, 
		output_MAC_12_30, output_MAC_12_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_13_0, output_MAC_13_1, output_MAC_13_2, output_MAC_13_3, output_MAC_13_4, output_MAC_13_5, output_MAC_13_6, output_MAC_13_7, output_MAC_13_8, output_MAC_13_9, 
		output_MAC_13_10, output_MAC_13_11, output_MAC_13_12, output_MAC_13_13, output_MAC_13_14, output_MAC_13_15, output_MAC_13_16, output_MAC_13_17, output_MAC_13_18, output_MAC_13_19, 
		output_MAC_13_20, output_MAC_13_21, output_MAC_13_22, output_MAC_13_23, output_MAC_13_24, output_MAC_13_25, output_MAC_13_26, output_MAC_13_27, output_MAC_13_28, output_MAC_13_29, 
		output_MAC_13_30, output_MAC_13_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_14_0, output_MAC_14_1, output_MAC_14_2, output_MAC_14_3, output_MAC_14_4, output_MAC_14_5, output_MAC_14_6, output_MAC_14_7, output_MAC_14_8, output_MAC_14_9, 
		output_MAC_14_10, output_MAC_14_11, output_MAC_14_12, output_MAC_14_13, output_MAC_14_14, output_MAC_14_15, output_MAC_14_16, output_MAC_14_17, output_MAC_14_18, output_MAC_14_19, 
		output_MAC_14_20, output_MAC_14_21, output_MAC_14_22, output_MAC_14_23, output_MAC_14_24, output_MAC_14_25, output_MAC_14_26, output_MAC_14_27, output_MAC_14_28, output_MAC_14_29, 
		output_MAC_14_30, output_MAC_14_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_15_0, output_MAC_15_1, output_MAC_15_2, output_MAC_15_3, output_MAC_15_4, output_MAC_15_5, output_MAC_15_6, output_MAC_15_7, output_MAC_15_8, output_MAC_15_9, 
		output_MAC_15_10, output_MAC_15_11, output_MAC_15_12, output_MAC_15_13, output_MAC_15_14, output_MAC_15_15, output_MAC_15_16, output_MAC_15_17, output_MAC_15_18, output_MAC_15_19, 
		output_MAC_15_20, output_MAC_15_21, output_MAC_15_22, output_MAC_15_23, output_MAC_15_24, output_MAC_15_25, output_MAC_15_26, output_MAC_15_27, output_MAC_15_28, output_MAC_15_29, 
		output_MAC_15_30, output_MAC_15_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_16_0, output_MAC_16_1, output_MAC_16_2, output_MAC_16_3, output_MAC_16_4, output_MAC_16_5, output_MAC_16_6, output_MAC_16_7, output_MAC_16_8, output_MAC_16_9, 
		output_MAC_16_10, output_MAC_16_11, output_MAC_16_12, output_MAC_16_13, output_MAC_16_14, output_MAC_16_15, output_MAC_16_16, output_MAC_16_17, output_MAC_16_18, output_MAC_16_19, 
		output_MAC_16_20, output_MAC_16_21, output_MAC_16_22, output_MAC_16_23, output_MAC_16_24, output_MAC_16_25, output_MAC_16_26, output_MAC_16_27, output_MAC_16_28, output_MAC_16_29, 
		output_MAC_16_30, output_MAC_16_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_17_0, output_MAC_17_1, output_MAC_17_2, output_MAC_17_3, output_MAC_17_4, output_MAC_17_5, output_MAC_17_6, output_MAC_17_7, output_MAC_17_8, output_MAC_17_9, 
		output_MAC_17_10, output_MAC_17_11, output_MAC_17_12, output_MAC_17_13, output_MAC_17_14, output_MAC_17_15, output_MAC_17_16, output_MAC_17_17, output_MAC_17_18, output_MAC_17_19, 
		output_MAC_17_20, output_MAC_17_21, output_MAC_17_22, output_MAC_17_23, output_MAC_17_24, output_MAC_17_25, output_MAC_17_26, output_MAC_17_27, output_MAC_17_28, output_MAC_17_29, 
		output_MAC_17_30, output_MAC_17_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_18_0, output_MAC_18_1, output_MAC_18_2, output_MAC_18_3, output_MAC_18_4, output_MAC_18_5, output_MAC_18_6, output_MAC_18_7, output_MAC_18_8, output_MAC_18_9, 
		output_MAC_18_10, output_MAC_18_11, output_MAC_18_12, output_MAC_18_13, output_MAC_18_14, output_MAC_18_15, output_MAC_18_16, output_MAC_18_17, output_MAC_18_18, output_MAC_18_19, 
		output_MAC_18_20, output_MAC_18_21, output_MAC_18_22, output_MAC_18_23, output_MAC_18_24, output_MAC_18_25, output_MAC_18_26, output_MAC_18_27, output_MAC_18_28, output_MAC_18_29, 
		output_MAC_18_30, output_MAC_18_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_19_0, output_MAC_19_1, output_MAC_19_2, output_MAC_19_3, output_MAC_19_4, output_MAC_19_5, output_MAC_19_6, output_MAC_19_7, output_MAC_19_8, output_MAC_19_9, 
		output_MAC_19_10, output_MAC_19_11, output_MAC_19_12, output_MAC_19_13, output_MAC_19_14, output_MAC_19_15, output_MAC_19_16, output_MAC_19_17, output_MAC_19_18, output_MAC_19_19, 
		output_MAC_19_20, output_MAC_19_21, output_MAC_19_22, output_MAC_19_23, output_MAC_19_24, output_MAC_19_25, output_MAC_19_26, output_MAC_19_27, output_MAC_19_28, output_MAC_19_29, 
		output_MAC_19_30, output_MAC_19_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_20_0, output_MAC_20_1, output_MAC_20_2, output_MAC_20_3, output_MAC_20_4, output_MAC_20_5, output_MAC_20_6, output_MAC_20_7, output_MAC_20_8, output_MAC_20_9, 
		output_MAC_20_10, output_MAC_20_11, output_MAC_20_12, output_MAC_20_13, output_MAC_20_14, output_MAC_20_15, output_MAC_20_16, output_MAC_20_17, output_MAC_20_18, output_MAC_20_19, 
		output_MAC_20_20, output_MAC_20_21, output_MAC_20_22, output_MAC_20_23, output_MAC_20_24, output_MAC_20_25, output_MAC_20_26, output_MAC_20_27, output_MAC_20_28, output_MAC_20_29, 
		output_MAC_20_30, output_MAC_20_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_21_0, output_MAC_21_1, output_MAC_21_2, output_MAC_21_3, output_MAC_21_4, output_MAC_21_5, output_MAC_21_6, output_MAC_21_7, output_MAC_21_8, output_MAC_21_9, 
		output_MAC_21_10, output_MAC_21_11, output_MAC_21_12, output_MAC_21_13, output_MAC_21_14, output_MAC_21_15, output_MAC_21_16, output_MAC_21_17, output_MAC_21_18, output_MAC_21_19, 
		output_MAC_21_20, output_MAC_21_21, output_MAC_21_22, output_MAC_21_23, output_MAC_21_24, output_MAC_21_25, output_MAC_21_26, output_MAC_21_27, output_MAC_21_28, output_MAC_21_29, 
		output_MAC_21_30, output_MAC_21_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_22_0, output_MAC_22_1, output_MAC_22_2, output_MAC_22_3, output_MAC_22_4, output_MAC_22_5, output_MAC_22_6, output_MAC_22_7, output_MAC_22_8, output_MAC_22_9, 
		output_MAC_22_10, output_MAC_22_11, output_MAC_22_12, output_MAC_22_13, output_MAC_22_14, output_MAC_22_15, output_MAC_22_16, output_MAC_22_17, output_MAC_22_18, output_MAC_22_19, 
		output_MAC_22_20, output_MAC_22_21, output_MAC_22_22, output_MAC_22_23, output_MAC_22_24, output_MAC_22_25, output_MAC_22_26, output_MAC_22_27, output_MAC_22_28, output_MAC_22_29, 
		output_MAC_22_30, output_MAC_22_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_23_0, output_MAC_23_1, output_MAC_23_2, output_MAC_23_3, output_MAC_23_4, output_MAC_23_5, output_MAC_23_6, output_MAC_23_7, output_MAC_23_8, output_MAC_23_9, 
		output_MAC_23_10, output_MAC_23_11, output_MAC_23_12, output_MAC_23_13, output_MAC_23_14, output_MAC_23_15, output_MAC_23_16, output_MAC_23_17, output_MAC_23_18, output_MAC_23_19, 
		output_MAC_23_20, output_MAC_23_21, output_MAC_23_22, output_MAC_23_23, output_MAC_23_24, output_MAC_23_25, output_MAC_23_26, output_MAC_23_27, output_MAC_23_28, output_MAC_23_29, 
		output_MAC_23_30, output_MAC_23_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_24_0, output_MAC_24_1, output_MAC_24_2, output_MAC_24_3, output_MAC_24_4, output_MAC_24_5, output_MAC_24_6, output_MAC_24_7, output_MAC_24_8, output_MAC_24_9, 
		output_MAC_24_10, output_MAC_24_11, output_MAC_24_12, output_MAC_24_13, output_MAC_24_14, output_MAC_24_15, output_MAC_24_16, output_MAC_24_17, output_MAC_24_18, output_MAC_24_19, 
		output_MAC_24_20, output_MAC_24_21, output_MAC_24_22, output_MAC_24_23, output_MAC_24_24, output_MAC_24_25, output_MAC_24_26, output_MAC_24_27, output_MAC_24_28, output_MAC_24_29, 
		output_MAC_24_30, output_MAC_24_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_25_0, output_MAC_25_1, output_MAC_25_2, output_MAC_25_3, output_MAC_25_4, output_MAC_25_5, output_MAC_25_6, output_MAC_25_7, output_MAC_25_8, output_MAC_25_9, 
		output_MAC_25_10, output_MAC_25_11, output_MAC_25_12, output_MAC_25_13, output_MAC_25_14, output_MAC_25_15, output_MAC_25_16, output_MAC_25_17, output_MAC_25_18, output_MAC_25_19, 
		output_MAC_25_20, output_MAC_25_21, output_MAC_25_22, output_MAC_25_23, output_MAC_25_24, output_MAC_25_25, output_MAC_25_26, output_MAC_25_27, output_MAC_25_28, output_MAC_25_29, 
		output_MAC_25_30, output_MAC_25_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_26_0, output_MAC_26_1, output_MAC_26_2, output_MAC_26_3, output_MAC_26_4, output_MAC_26_5, output_MAC_26_6, output_MAC_26_7, output_MAC_26_8, output_MAC_26_9, 
		output_MAC_26_10, output_MAC_26_11, output_MAC_26_12, output_MAC_26_13, output_MAC_26_14, output_MAC_26_15, output_MAC_26_16, output_MAC_26_17, output_MAC_26_18, output_MAC_26_19, 
		output_MAC_26_20, output_MAC_26_21, output_MAC_26_22, output_MAC_26_23, output_MAC_26_24, output_MAC_26_25, output_MAC_26_26, output_MAC_26_27, output_MAC_26_28, output_MAC_26_29, 
		output_MAC_26_30, output_MAC_26_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_27_0, output_MAC_27_1, output_MAC_27_2, output_MAC_27_3, output_MAC_27_4, output_MAC_27_5, output_MAC_27_6, output_MAC_27_7, output_MAC_27_8, output_MAC_27_9, 
		output_MAC_27_10, output_MAC_27_11, output_MAC_27_12, output_MAC_27_13, output_MAC_27_14, output_MAC_27_15, output_MAC_27_16, output_MAC_27_17, output_MAC_27_18, output_MAC_27_19, 
		output_MAC_27_20, output_MAC_27_21, output_MAC_27_22, output_MAC_27_23, output_MAC_27_24, output_MAC_27_25, output_MAC_27_26, output_MAC_27_27, output_MAC_27_28, output_MAC_27_29, 
		output_MAC_27_30, output_MAC_27_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_28_0, output_MAC_28_1, output_MAC_28_2, output_MAC_28_3, output_MAC_28_4, output_MAC_28_5, output_MAC_28_6, output_MAC_28_7, output_MAC_28_8, output_MAC_28_9, 
		output_MAC_28_10, output_MAC_28_11, output_MAC_28_12, output_MAC_28_13, output_MAC_28_14, output_MAC_28_15, output_MAC_28_16, output_MAC_28_17, output_MAC_28_18, output_MAC_28_19, 
		output_MAC_28_20, output_MAC_28_21, output_MAC_28_22, output_MAC_28_23, output_MAC_28_24, output_MAC_28_25, output_MAC_28_26, output_MAC_28_27, output_MAC_28_28, output_MAC_28_29, 
		output_MAC_28_30, output_MAC_28_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_29_0, output_MAC_29_1, output_MAC_29_2, output_MAC_29_3, output_MAC_29_4, output_MAC_29_5, output_MAC_29_6, output_MAC_29_7, output_MAC_29_8, output_MAC_29_9, 
		output_MAC_29_10, output_MAC_29_11, output_MAC_29_12, output_MAC_29_13, output_MAC_29_14, output_MAC_29_15, output_MAC_29_16, output_MAC_29_17, output_MAC_29_18, output_MAC_29_19, 
		output_MAC_29_20, output_MAC_29_21, output_MAC_29_22, output_MAC_29_23, output_MAC_29_24, output_MAC_29_25, output_MAC_29_26, output_MAC_29_27, output_MAC_29_28, output_MAC_29_29, 
		output_MAC_29_30, output_MAC_29_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_30_0, output_MAC_30_1, output_MAC_30_2, output_MAC_30_3, output_MAC_30_4, output_MAC_30_5, output_MAC_30_6, output_MAC_30_7, output_MAC_30_8, output_MAC_30_9, 
		output_MAC_30_10, output_MAC_30_11, output_MAC_30_12, output_MAC_30_13, output_MAC_30_14, output_MAC_30_15, output_MAC_30_16, output_MAC_30_17, output_MAC_30_18, output_MAC_30_19, 
		output_MAC_30_20, output_MAC_30_21, output_MAC_30_22, output_MAC_30_23, output_MAC_30_24, output_MAC_30_25, output_MAC_30_26, output_MAC_30_27, output_MAC_30_28, output_MAC_30_29, 
		output_MAC_30_30, output_MAC_30_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_31_0, output_MAC_31_1, output_MAC_31_2, output_MAC_31_3, output_MAC_31_4, output_MAC_31_5, output_MAC_31_6, output_MAC_31_7, output_MAC_31_8, output_MAC_31_9, 
		output_MAC_31_10, output_MAC_31_11, output_MAC_31_12, output_MAC_31_13, output_MAC_31_14, output_MAC_31_15, output_MAC_31_16, output_MAC_31_17, output_MAC_31_18, output_MAC_31_19, 
		output_MAC_31_20, output_MAC_31_21, output_MAC_31_22, output_MAC_31_23, output_MAC_31_24, output_MAC_31_25, output_MAC_31_26, output_MAC_31_27, output_MAC_31_28, output_MAC_31_29, 
		output_MAC_31_30, output_MAC_31_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_32_0, output_MAC_32_1, output_MAC_32_2, output_MAC_32_3, output_MAC_32_4, output_MAC_32_5, output_MAC_32_6, output_MAC_32_7, output_MAC_32_8, output_MAC_32_9, 
		output_MAC_32_10, output_MAC_32_11, output_MAC_32_12, output_MAC_32_13, output_MAC_32_14, output_MAC_32_15, output_MAC_32_16, output_MAC_32_17, output_MAC_32_18, output_MAC_32_19, 
		output_MAC_32_20, output_MAC_32_21, output_MAC_32_22, output_MAC_32_23, output_MAC_32_24, output_MAC_32_25, output_MAC_32_26, output_MAC_32_27, output_MAC_32_28, output_MAC_32_29, 
		output_MAC_32_30, output_MAC_32_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_33_0, output_MAC_33_1, output_MAC_33_2, output_MAC_33_3, output_MAC_33_4, output_MAC_33_5, output_MAC_33_6, output_MAC_33_7, output_MAC_33_8, output_MAC_33_9, 
		output_MAC_33_10, output_MAC_33_11, output_MAC_33_12, output_MAC_33_13, output_MAC_33_14, output_MAC_33_15, output_MAC_33_16, output_MAC_33_17, output_MAC_33_18, output_MAC_33_19, 
		output_MAC_33_20, output_MAC_33_21, output_MAC_33_22, output_MAC_33_23, output_MAC_33_24, output_MAC_33_25, output_MAC_33_26, output_MAC_33_27, output_MAC_33_28, output_MAC_33_29, 
		output_MAC_33_30, output_MAC_33_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_34_0, output_MAC_34_1, output_MAC_34_2, output_MAC_34_3, output_MAC_34_4, output_MAC_34_5, output_MAC_34_6, output_MAC_34_7, output_MAC_34_8, output_MAC_34_9, 
		output_MAC_34_10, output_MAC_34_11, output_MAC_34_12, output_MAC_34_13, output_MAC_34_14, output_MAC_34_15, output_MAC_34_16, output_MAC_34_17, output_MAC_34_18, output_MAC_34_19, 
		output_MAC_34_20, output_MAC_34_21, output_MAC_34_22, output_MAC_34_23, output_MAC_34_24, output_MAC_34_25, output_MAC_34_26, output_MAC_34_27, output_MAC_34_28, output_MAC_34_29, 
		output_MAC_34_30, output_MAC_34_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_35_0, output_MAC_35_1, output_MAC_35_2, output_MAC_35_3, output_MAC_35_4, output_MAC_35_5, output_MAC_35_6, output_MAC_35_7, output_MAC_35_8, output_MAC_35_9, 
		output_MAC_35_10, output_MAC_35_11, output_MAC_35_12, output_MAC_35_13, output_MAC_35_14, output_MAC_35_15, output_MAC_35_16, output_MAC_35_17, output_MAC_35_18, output_MAC_35_19, 
		output_MAC_35_20, output_MAC_35_21, output_MAC_35_22, output_MAC_35_23, output_MAC_35_24, output_MAC_35_25, output_MAC_35_26, output_MAC_35_27, output_MAC_35_28, output_MAC_35_29, 
		output_MAC_35_30, output_MAC_35_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_36_0, output_MAC_36_1, output_MAC_36_2, output_MAC_36_3, output_MAC_36_4, output_MAC_36_5, output_MAC_36_6, output_MAC_36_7, output_MAC_36_8, output_MAC_36_9, 
		output_MAC_36_10, output_MAC_36_11, output_MAC_36_12, output_MAC_36_13, output_MAC_36_14, output_MAC_36_15, output_MAC_36_16, output_MAC_36_17, output_MAC_36_18, output_MAC_36_19, 
		output_MAC_36_20, output_MAC_36_21, output_MAC_36_22, output_MAC_36_23, output_MAC_36_24, output_MAC_36_25, output_MAC_36_26, output_MAC_36_27, output_MAC_36_28, output_MAC_36_29, 
		output_MAC_36_30, output_MAC_36_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_37_0, output_MAC_37_1, output_MAC_37_2, output_MAC_37_3, output_MAC_37_4, output_MAC_37_5, output_MAC_37_6, output_MAC_37_7, output_MAC_37_8, output_MAC_37_9, 
		output_MAC_37_10, output_MAC_37_11, output_MAC_37_12, output_MAC_37_13, output_MAC_37_14, output_MAC_37_15, output_MAC_37_16, output_MAC_37_17, output_MAC_37_18, output_MAC_37_19, 
		output_MAC_37_20, output_MAC_37_21, output_MAC_37_22, output_MAC_37_23, output_MAC_37_24, output_MAC_37_25, output_MAC_37_26, output_MAC_37_27, output_MAC_37_28, output_MAC_37_29, 
		output_MAC_37_30, output_MAC_37_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_38_0, output_MAC_38_1, output_MAC_38_2, output_MAC_38_3, output_MAC_38_4, output_MAC_38_5, output_MAC_38_6, output_MAC_38_7, output_MAC_38_8, output_MAC_38_9, 
		output_MAC_38_10, output_MAC_38_11, output_MAC_38_12, output_MAC_38_13, output_MAC_38_14, output_MAC_38_15, output_MAC_38_16, output_MAC_38_17, output_MAC_38_18, output_MAC_38_19, 
		output_MAC_38_20, output_MAC_38_21, output_MAC_38_22, output_MAC_38_23, output_MAC_38_24, output_MAC_38_25, output_MAC_38_26, output_MAC_38_27, output_MAC_38_28, output_MAC_38_29, 
		output_MAC_38_30, output_MAC_38_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_39_0, output_MAC_39_1, output_MAC_39_2, output_MAC_39_3, output_MAC_39_4, output_MAC_39_5, output_MAC_39_6, output_MAC_39_7, output_MAC_39_8, output_MAC_39_9, 
		output_MAC_39_10, output_MAC_39_11, output_MAC_39_12, output_MAC_39_13, output_MAC_39_14, output_MAC_39_15, output_MAC_39_16, output_MAC_39_17, output_MAC_39_18, output_MAC_39_19, 
		output_MAC_39_20, output_MAC_39_21, output_MAC_39_22, output_MAC_39_23, output_MAC_39_24, output_MAC_39_25, output_MAC_39_26, output_MAC_39_27, output_MAC_39_28, output_MAC_39_29, 
		output_MAC_39_30, output_MAC_39_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_40_0, output_MAC_40_1, output_MAC_40_2, output_MAC_40_3, output_MAC_40_4, output_MAC_40_5, output_MAC_40_6, output_MAC_40_7, output_MAC_40_8, output_MAC_40_9, 
		output_MAC_40_10, output_MAC_40_11, output_MAC_40_12, output_MAC_40_13, output_MAC_40_14, output_MAC_40_15, output_MAC_40_16, output_MAC_40_17, output_MAC_40_18, output_MAC_40_19, 
		output_MAC_40_20, output_MAC_40_21, output_MAC_40_22, output_MAC_40_23, output_MAC_40_24, output_MAC_40_25, output_MAC_40_26, output_MAC_40_27, output_MAC_40_28, output_MAC_40_29, 
		output_MAC_40_30, output_MAC_40_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_41_0, output_MAC_41_1, output_MAC_41_2, output_MAC_41_3, output_MAC_41_4, output_MAC_41_5, output_MAC_41_6, output_MAC_41_7, output_MAC_41_8, output_MAC_41_9, 
		output_MAC_41_10, output_MAC_41_11, output_MAC_41_12, output_MAC_41_13, output_MAC_41_14, output_MAC_41_15, output_MAC_41_16, output_MAC_41_17, output_MAC_41_18, output_MAC_41_19, 
		output_MAC_41_20, output_MAC_41_21, output_MAC_41_22, output_MAC_41_23, output_MAC_41_24, output_MAC_41_25, output_MAC_41_26, output_MAC_41_27, output_MAC_41_28, output_MAC_41_29, 
		output_MAC_41_30, output_MAC_41_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_42_0, output_MAC_42_1, output_MAC_42_2, output_MAC_42_3, output_MAC_42_4, output_MAC_42_5, output_MAC_42_6, output_MAC_42_7, output_MAC_42_8, output_MAC_42_9, 
		output_MAC_42_10, output_MAC_42_11, output_MAC_42_12, output_MAC_42_13, output_MAC_42_14, output_MAC_42_15, output_MAC_42_16, output_MAC_42_17, output_MAC_42_18, output_MAC_42_19, 
		output_MAC_42_20, output_MAC_42_21, output_MAC_42_22, output_MAC_42_23, output_MAC_42_24, output_MAC_42_25, output_MAC_42_26, output_MAC_42_27, output_MAC_42_28, output_MAC_42_29, 
		output_MAC_42_30, output_MAC_42_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_43_0, output_MAC_43_1, output_MAC_43_2, output_MAC_43_3, output_MAC_43_4, output_MAC_43_5, output_MAC_43_6, output_MAC_43_7, output_MAC_43_8, output_MAC_43_9, 
		output_MAC_43_10, output_MAC_43_11, output_MAC_43_12, output_MAC_43_13, output_MAC_43_14, output_MAC_43_15, output_MAC_43_16, output_MAC_43_17, output_MAC_43_18, output_MAC_43_19, 
		output_MAC_43_20, output_MAC_43_21, output_MAC_43_22, output_MAC_43_23, output_MAC_43_24, output_MAC_43_25, output_MAC_43_26, output_MAC_43_27, output_MAC_43_28, output_MAC_43_29, 
		output_MAC_43_30, output_MAC_43_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_44_0, output_MAC_44_1, output_MAC_44_2, output_MAC_44_3, output_MAC_44_4, output_MAC_44_5, output_MAC_44_6, output_MAC_44_7, output_MAC_44_8, output_MAC_44_9, 
		output_MAC_44_10, output_MAC_44_11, output_MAC_44_12, output_MAC_44_13, output_MAC_44_14, output_MAC_44_15, output_MAC_44_16, output_MAC_44_17, output_MAC_44_18, output_MAC_44_19, 
		output_MAC_44_20, output_MAC_44_21, output_MAC_44_22, output_MAC_44_23, output_MAC_44_24, output_MAC_44_25, output_MAC_44_26, output_MAC_44_27, output_MAC_44_28, output_MAC_44_29, 
		output_MAC_44_30, output_MAC_44_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_45_0, output_MAC_45_1, output_MAC_45_2, output_MAC_45_3, output_MAC_45_4, output_MAC_45_5, output_MAC_45_6, output_MAC_45_7, output_MAC_45_8, output_MAC_45_9, 
		output_MAC_45_10, output_MAC_45_11, output_MAC_45_12, output_MAC_45_13, output_MAC_45_14, output_MAC_45_15, output_MAC_45_16, output_MAC_45_17, output_MAC_45_18, output_MAC_45_19, 
		output_MAC_45_20, output_MAC_45_21, output_MAC_45_22, output_MAC_45_23, output_MAC_45_24, output_MAC_45_25, output_MAC_45_26, output_MAC_45_27, output_MAC_45_28, output_MAC_45_29, 
		output_MAC_45_30, output_MAC_45_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_46_0, output_MAC_46_1, output_MAC_46_2, output_MAC_46_3, output_MAC_46_4, output_MAC_46_5, output_MAC_46_6, output_MAC_46_7, output_MAC_46_8, output_MAC_46_9, 
		output_MAC_46_10, output_MAC_46_11, output_MAC_46_12, output_MAC_46_13, output_MAC_46_14, output_MAC_46_15, output_MAC_46_16, output_MAC_46_17, output_MAC_46_18, output_MAC_46_19, 
		output_MAC_46_20, output_MAC_46_21, output_MAC_46_22, output_MAC_46_23, output_MAC_46_24, output_MAC_46_25, output_MAC_46_26, output_MAC_46_27, output_MAC_46_28, output_MAC_46_29, 
		output_MAC_46_30, output_MAC_46_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_47_0, output_MAC_47_1, output_MAC_47_2, output_MAC_47_3, output_MAC_47_4, output_MAC_47_5, output_MAC_47_6, output_MAC_47_7, output_MAC_47_8, output_MAC_47_9, 
		output_MAC_47_10, output_MAC_47_11, output_MAC_47_12, output_MAC_47_13, output_MAC_47_14, output_MAC_47_15, output_MAC_47_16, output_MAC_47_17, output_MAC_47_18, output_MAC_47_19, 
		output_MAC_47_20, output_MAC_47_21, output_MAC_47_22, output_MAC_47_23, output_MAC_47_24, output_MAC_47_25, output_MAC_47_26, output_MAC_47_27, output_MAC_47_28, output_MAC_47_29, 
		output_MAC_47_30, output_MAC_47_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_48_0, output_MAC_48_1, output_MAC_48_2, output_MAC_48_3, output_MAC_48_4, output_MAC_48_5, output_MAC_48_6, output_MAC_48_7, output_MAC_48_8, output_MAC_48_9, 
		output_MAC_48_10, output_MAC_48_11, output_MAC_48_12, output_MAC_48_13, output_MAC_48_14, output_MAC_48_15, output_MAC_48_16, output_MAC_48_17, output_MAC_48_18, output_MAC_48_19, 
		output_MAC_48_20, output_MAC_48_21, output_MAC_48_22, output_MAC_48_23, output_MAC_48_24, output_MAC_48_25, output_MAC_48_26, output_MAC_48_27, output_MAC_48_28, output_MAC_48_29, 
		output_MAC_48_30, output_MAC_48_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_49_0, output_MAC_49_1, output_MAC_49_2, output_MAC_49_3, output_MAC_49_4, output_MAC_49_5, output_MAC_49_6, output_MAC_49_7, output_MAC_49_8, output_MAC_49_9, 
		output_MAC_49_10, output_MAC_49_11, output_MAC_49_12, output_MAC_49_13, output_MAC_49_14, output_MAC_49_15, output_MAC_49_16, output_MAC_49_17, output_MAC_49_18, output_MAC_49_19, 
		output_MAC_49_20, output_MAC_49_21, output_MAC_49_22, output_MAC_49_23, output_MAC_49_24, output_MAC_49_25, output_MAC_49_26, output_MAC_49_27, output_MAC_49_28, output_MAC_49_29, 
		output_MAC_49_30, output_MAC_49_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_50_0, output_MAC_50_1, output_MAC_50_2, output_MAC_50_3, output_MAC_50_4, output_MAC_50_5, output_MAC_50_6, output_MAC_50_7, output_MAC_50_8, output_MAC_50_9, 
		output_MAC_50_10, output_MAC_50_11, output_MAC_50_12, output_MAC_50_13, output_MAC_50_14, output_MAC_50_15, output_MAC_50_16, output_MAC_50_17, output_MAC_50_18, output_MAC_50_19, 
		output_MAC_50_20, output_MAC_50_21, output_MAC_50_22, output_MAC_50_23, output_MAC_50_24, output_MAC_50_25, output_MAC_50_26, output_MAC_50_27, output_MAC_50_28, output_MAC_50_29, 
		output_MAC_50_30, output_MAC_50_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_51_0, output_MAC_51_1, output_MAC_51_2, output_MAC_51_3, output_MAC_51_4, output_MAC_51_5, output_MAC_51_6, output_MAC_51_7, output_MAC_51_8, output_MAC_51_9, 
		output_MAC_51_10, output_MAC_51_11, output_MAC_51_12, output_MAC_51_13, output_MAC_51_14, output_MAC_51_15, output_MAC_51_16, output_MAC_51_17, output_MAC_51_18, output_MAC_51_19, 
		output_MAC_51_20, output_MAC_51_21, output_MAC_51_22, output_MAC_51_23, output_MAC_51_24, output_MAC_51_25, output_MAC_51_26, output_MAC_51_27, output_MAC_51_28, output_MAC_51_29, 
		output_MAC_51_30, output_MAC_51_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_52_0, output_MAC_52_1, output_MAC_52_2, output_MAC_52_3, output_MAC_52_4, output_MAC_52_5, output_MAC_52_6, output_MAC_52_7, output_MAC_52_8, output_MAC_52_9, 
		output_MAC_52_10, output_MAC_52_11, output_MAC_52_12, output_MAC_52_13, output_MAC_52_14, output_MAC_52_15, output_MAC_52_16, output_MAC_52_17, output_MAC_52_18, output_MAC_52_19, 
		output_MAC_52_20, output_MAC_52_21, output_MAC_52_22, output_MAC_52_23, output_MAC_52_24, output_MAC_52_25, output_MAC_52_26, output_MAC_52_27, output_MAC_52_28, output_MAC_52_29, 
		output_MAC_52_30, output_MAC_52_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_53_0, output_MAC_53_1, output_MAC_53_2, output_MAC_53_3, output_MAC_53_4, output_MAC_53_5, output_MAC_53_6, output_MAC_53_7, output_MAC_53_8, output_MAC_53_9, 
		output_MAC_53_10, output_MAC_53_11, output_MAC_53_12, output_MAC_53_13, output_MAC_53_14, output_MAC_53_15, output_MAC_53_16, output_MAC_53_17, output_MAC_53_18, output_MAC_53_19, 
		output_MAC_53_20, output_MAC_53_21, output_MAC_53_22, output_MAC_53_23, output_MAC_53_24, output_MAC_53_25, output_MAC_53_26, output_MAC_53_27, output_MAC_53_28, output_MAC_53_29, 
		output_MAC_53_30, output_MAC_53_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_54_0, output_MAC_54_1, output_MAC_54_2, output_MAC_54_3, output_MAC_54_4, output_MAC_54_5, output_MAC_54_6, output_MAC_54_7, output_MAC_54_8, output_MAC_54_9, 
		output_MAC_54_10, output_MAC_54_11, output_MAC_54_12, output_MAC_54_13, output_MAC_54_14, output_MAC_54_15, output_MAC_54_16, output_MAC_54_17, output_MAC_54_18, output_MAC_54_19, 
		output_MAC_54_20, output_MAC_54_21, output_MAC_54_22, output_MAC_54_23, output_MAC_54_24, output_MAC_54_25, output_MAC_54_26, output_MAC_54_27, output_MAC_54_28, output_MAC_54_29, 
		output_MAC_54_30, output_MAC_54_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_55_0, output_MAC_55_1, output_MAC_55_2, output_MAC_55_3, output_MAC_55_4, output_MAC_55_5, output_MAC_55_6, output_MAC_55_7, output_MAC_55_8, output_MAC_55_9, 
		output_MAC_55_10, output_MAC_55_11, output_MAC_55_12, output_MAC_55_13, output_MAC_55_14, output_MAC_55_15, output_MAC_55_16, output_MAC_55_17, output_MAC_55_18, output_MAC_55_19, 
		output_MAC_55_20, output_MAC_55_21, output_MAC_55_22, output_MAC_55_23, output_MAC_55_24, output_MAC_55_25, output_MAC_55_26, output_MAC_55_27, output_MAC_55_28, output_MAC_55_29, 
		output_MAC_55_30, output_MAC_55_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_56_0, output_MAC_56_1, output_MAC_56_2, output_MAC_56_3, output_MAC_56_4, output_MAC_56_5, output_MAC_56_6, output_MAC_56_7, output_MAC_56_8, output_MAC_56_9, 
		output_MAC_56_10, output_MAC_56_11, output_MAC_56_12, output_MAC_56_13, output_MAC_56_14, output_MAC_56_15, output_MAC_56_16, output_MAC_56_17, output_MAC_56_18, output_MAC_56_19, 
		output_MAC_56_20, output_MAC_56_21, output_MAC_56_22, output_MAC_56_23, output_MAC_56_24, output_MAC_56_25, output_MAC_56_26, output_MAC_56_27, output_MAC_56_28, output_MAC_56_29, 
		output_MAC_56_30, output_MAC_56_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_57_0, output_MAC_57_1, output_MAC_57_2, output_MAC_57_3, output_MAC_57_4, output_MAC_57_5, output_MAC_57_6, output_MAC_57_7, output_MAC_57_8, output_MAC_57_9, 
		output_MAC_57_10, output_MAC_57_11, output_MAC_57_12, output_MAC_57_13, output_MAC_57_14, output_MAC_57_15, output_MAC_57_16, output_MAC_57_17, output_MAC_57_18, output_MAC_57_19, 
		output_MAC_57_20, output_MAC_57_21, output_MAC_57_22, output_MAC_57_23, output_MAC_57_24, output_MAC_57_25, output_MAC_57_26, output_MAC_57_27, output_MAC_57_28, output_MAC_57_29, 
		output_MAC_57_30, output_MAC_57_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_58_0, output_MAC_58_1, output_MAC_58_2, output_MAC_58_3, output_MAC_58_4, output_MAC_58_5, output_MAC_58_6, output_MAC_58_7, output_MAC_58_8, output_MAC_58_9, 
		output_MAC_58_10, output_MAC_58_11, output_MAC_58_12, output_MAC_58_13, output_MAC_58_14, output_MAC_58_15, output_MAC_58_16, output_MAC_58_17, output_MAC_58_18, output_MAC_58_19, 
		output_MAC_58_20, output_MAC_58_21, output_MAC_58_22, output_MAC_58_23, output_MAC_58_24, output_MAC_58_25, output_MAC_58_26, output_MAC_58_27, output_MAC_58_28, output_MAC_58_29, 
		output_MAC_58_30, output_MAC_58_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_59_0, output_MAC_59_1, output_MAC_59_2, output_MAC_59_3, output_MAC_59_4, output_MAC_59_5, output_MAC_59_6, output_MAC_59_7, output_MAC_59_8, output_MAC_59_9, 
		output_MAC_59_10, output_MAC_59_11, output_MAC_59_12, output_MAC_59_13, output_MAC_59_14, output_MAC_59_15, output_MAC_59_16, output_MAC_59_17, output_MAC_59_18, output_MAC_59_19, 
		output_MAC_59_20, output_MAC_59_21, output_MAC_59_22, output_MAC_59_23, output_MAC_59_24, output_MAC_59_25, output_MAC_59_26, output_MAC_59_27, output_MAC_59_28, output_MAC_59_29, 
		output_MAC_59_30, output_MAC_59_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_60_0, output_MAC_60_1, output_MAC_60_2, output_MAC_60_3, output_MAC_60_4, output_MAC_60_5, output_MAC_60_6, output_MAC_60_7, output_MAC_60_8, output_MAC_60_9, 
		output_MAC_60_10, output_MAC_60_11, output_MAC_60_12, output_MAC_60_13, output_MAC_60_14, output_MAC_60_15, output_MAC_60_16, output_MAC_60_17, output_MAC_60_18, output_MAC_60_19, 
		output_MAC_60_20, output_MAC_60_21, output_MAC_60_22, output_MAC_60_23, output_MAC_60_24, output_MAC_60_25, output_MAC_60_26, output_MAC_60_27, output_MAC_60_28, output_MAC_60_29, 
		output_MAC_60_30, output_MAC_60_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_61_0, output_MAC_61_1, output_MAC_61_2, output_MAC_61_3, output_MAC_61_4, output_MAC_61_5, output_MAC_61_6, output_MAC_61_7, output_MAC_61_8, output_MAC_61_9, 
		output_MAC_61_10, output_MAC_61_11, output_MAC_61_12, output_MAC_61_13, output_MAC_61_14, output_MAC_61_15, output_MAC_61_16, output_MAC_61_17, output_MAC_61_18, output_MAC_61_19, 
		output_MAC_61_20, output_MAC_61_21, output_MAC_61_22, output_MAC_61_23, output_MAC_61_24, output_MAC_61_25, output_MAC_61_26, output_MAC_61_27, output_MAC_61_28, output_MAC_61_29, 
		output_MAC_61_30, output_MAC_61_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_62_0, output_MAC_62_1, output_MAC_62_2, output_MAC_62_3, output_MAC_62_4, output_MAC_62_5, output_MAC_62_6, output_MAC_62_7, output_MAC_62_8, output_MAC_62_9, 
		output_MAC_62_10, output_MAC_62_11, output_MAC_62_12, output_MAC_62_13, output_MAC_62_14, output_MAC_62_15, output_MAC_62_16, output_MAC_62_17, output_MAC_62_18, output_MAC_62_19, 
		output_MAC_62_20, output_MAC_62_21, output_MAC_62_22, output_MAC_62_23, output_MAC_62_24, output_MAC_62_25, output_MAC_62_26, output_MAC_62_27, output_MAC_62_28, output_MAC_62_29, 
		output_MAC_62_30, output_MAC_62_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_63_0, output_MAC_63_1, output_MAC_63_2, output_MAC_63_3, output_MAC_63_4, output_MAC_63_5, output_MAC_63_6, output_MAC_63_7, output_MAC_63_8, output_MAC_63_9, 
		output_MAC_63_10, output_MAC_63_11, output_MAC_63_12, output_MAC_63_13, output_MAC_63_14, output_MAC_63_15, output_MAC_63_16, output_MAC_63_17, output_MAC_63_18, output_MAC_63_19, 
		output_MAC_63_20, output_MAC_63_21, output_MAC_63_22, output_MAC_63_23, output_MAC_63_24, output_MAC_63_25, output_MAC_63_26, output_MAC_63_27, output_MAC_63_28, output_MAC_63_29, 
		output_MAC_63_30, output_MAC_63_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_64_0, output_MAC_64_1, output_MAC_64_2, output_MAC_64_3, output_MAC_64_4, output_MAC_64_5, output_MAC_64_6, output_MAC_64_7, output_MAC_64_8, output_MAC_64_9, 
		output_MAC_64_10, output_MAC_64_11, output_MAC_64_12, output_MAC_64_13, output_MAC_64_14, output_MAC_64_15, output_MAC_64_16, output_MAC_64_17, output_MAC_64_18, output_MAC_64_19, 
		output_MAC_64_20, output_MAC_64_21, output_MAC_64_22, output_MAC_64_23, output_MAC_64_24, output_MAC_64_25, output_MAC_64_26, output_MAC_64_27, output_MAC_64_28, output_MAC_64_29, 
		output_MAC_64_30, output_MAC_64_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_65_0, output_MAC_65_1, output_MAC_65_2, output_MAC_65_3, output_MAC_65_4, output_MAC_65_5, output_MAC_65_6, output_MAC_65_7, output_MAC_65_8, output_MAC_65_9, 
		output_MAC_65_10, output_MAC_65_11, output_MAC_65_12, output_MAC_65_13, output_MAC_65_14, output_MAC_65_15, output_MAC_65_16, output_MAC_65_17, output_MAC_65_18, output_MAC_65_19, 
		output_MAC_65_20, output_MAC_65_21, output_MAC_65_22, output_MAC_65_23, output_MAC_65_24, output_MAC_65_25, output_MAC_65_26, output_MAC_65_27, output_MAC_65_28, output_MAC_65_29, 
		output_MAC_65_30, output_MAC_65_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_66_0, output_MAC_66_1, output_MAC_66_2, output_MAC_66_3, output_MAC_66_4, output_MAC_66_5, output_MAC_66_6, output_MAC_66_7, output_MAC_66_8, output_MAC_66_9, 
		output_MAC_66_10, output_MAC_66_11, output_MAC_66_12, output_MAC_66_13, output_MAC_66_14, output_MAC_66_15, output_MAC_66_16, output_MAC_66_17, output_MAC_66_18, output_MAC_66_19, 
		output_MAC_66_20, output_MAC_66_21, output_MAC_66_22, output_MAC_66_23, output_MAC_66_24, output_MAC_66_25, output_MAC_66_26, output_MAC_66_27, output_MAC_66_28, output_MAC_66_29, 
		output_MAC_66_30, output_MAC_66_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_67_0, output_MAC_67_1, output_MAC_67_2, output_MAC_67_3, output_MAC_67_4, output_MAC_67_5, output_MAC_67_6, output_MAC_67_7, output_MAC_67_8, output_MAC_67_9, 
		output_MAC_67_10, output_MAC_67_11, output_MAC_67_12, output_MAC_67_13, output_MAC_67_14, output_MAC_67_15, output_MAC_67_16, output_MAC_67_17, output_MAC_67_18, output_MAC_67_19, 
		output_MAC_67_20, output_MAC_67_21, output_MAC_67_22, output_MAC_67_23, output_MAC_67_24, output_MAC_67_25, output_MAC_67_26, output_MAC_67_27, output_MAC_67_28, output_MAC_67_29, 
		output_MAC_67_30, output_MAC_67_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_68_0, output_MAC_68_1, output_MAC_68_2, output_MAC_68_3, output_MAC_68_4, output_MAC_68_5, output_MAC_68_6, output_MAC_68_7, output_MAC_68_8, output_MAC_68_9, 
		output_MAC_68_10, output_MAC_68_11, output_MAC_68_12, output_MAC_68_13, output_MAC_68_14, output_MAC_68_15, output_MAC_68_16, output_MAC_68_17, output_MAC_68_18, output_MAC_68_19, 
		output_MAC_68_20, output_MAC_68_21, output_MAC_68_22, output_MAC_68_23, output_MAC_68_24, output_MAC_68_25, output_MAC_68_26, output_MAC_68_27, output_MAC_68_28, output_MAC_68_29, 
		output_MAC_68_30, output_MAC_68_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_69_0, output_MAC_69_1, output_MAC_69_2, output_MAC_69_3, output_MAC_69_4, output_MAC_69_5, output_MAC_69_6, output_MAC_69_7, output_MAC_69_8, output_MAC_69_9, 
		output_MAC_69_10, output_MAC_69_11, output_MAC_69_12, output_MAC_69_13, output_MAC_69_14, output_MAC_69_15, output_MAC_69_16, output_MAC_69_17, output_MAC_69_18, output_MAC_69_19, 
		output_MAC_69_20, output_MAC_69_21, output_MAC_69_22, output_MAC_69_23, output_MAC_69_24, output_MAC_69_25, output_MAC_69_26, output_MAC_69_27, output_MAC_69_28, output_MAC_69_29, 
		output_MAC_69_30, output_MAC_69_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_70_0, output_MAC_70_1, output_MAC_70_2, output_MAC_70_3, output_MAC_70_4, output_MAC_70_5, output_MAC_70_6, output_MAC_70_7, output_MAC_70_8, output_MAC_70_9, 
		output_MAC_70_10, output_MAC_70_11, output_MAC_70_12, output_MAC_70_13, output_MAC_70_14, output_MAC_70_15, output_MAC_70_16, output_MAC_70_17, output_MAC_70_18, output_MAC_70_19, 
		output_MAC_70_20, output_MAC_70_21, output_MAC_70_22, output_MAC_70_23, output_MAC_70_24, output_MAC_70_25, output_MAC_70_26, output_MAC_70_27, output_MAC_70_28, output_MAC_70_29, 
		output_MAC_70_30, output_MAC_70_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_71_0, output_MAC_71_1, output_MAC_71_2, output_MAC_71_3, output_MAC_71_4, output_MAC_71_5, output_MAC_71_6, output_MAC_71_7, output_MAC_71_8, output_MAC_71_9, 
		output_MAC_71_10, output_MAC_71_11, output_MAC_71_12, output_MAC_71_13, output_MAC_71_14, output_MAC_71_15, output_MAC_71_16, output_MAC_71_17, output_MAC_71_18, output_MAC_71_19, 
		output_MAC_71_20, output_MAC_71_21, output_MAC_71_22, output_MAC_71_23, output_MAC_71_24, output_MAC_71_25, output_MAC_71_26, output_MAC_71_27, output_MAC_71_28, output_MAC_71_29, 
		output_MAC_71_30, output_MAC_71_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_72_0, output_MAC_72_1, output_MAC_72_2, output_MAC_72_3, output_MAC_72_4, output_MAC_72_5, output_MAC_72_6, output_MAC_72_7, output_MAC_72_8, output_MAC_72_9, 
		output_MAC_72_10, output_MAC_72_11, output_MAC_72_12, output_MAC_72_13, output_MAC_72_14, output_MAC_72_15, output_MAC_72_16, output_MAC_72_17, output_MAC_72_18, output_MAC_72_19, 
		output_MAC_72_20, output_MAC_72_21, output_MAC_72_22, output_MAC_72_23, output_MAC_72_24, output_MAC_72_25, output_MAC_72_26, output_MAC_72_27, output_MAC_72_28, output_MAC_72_29, 
		output_MAC_72_30, output_MAC_72_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_73_0, output_MAC_73_1, output_MAC_73_2, output_MAC_73_3, output_MAC_73_4, output_MAC_73_5, output_MAC_73_6, output_MAC_73_7, output_MAC_73_8, output_MAC_73_9, 
		output_MAC_73_10, output_MAC_73_11, output_MAC_73_12, output_MAC_73_13, output_MAC_73_14, output_MAC_73_15, output_MAC_73_16, output_MAC_73_17, output_MAC_73_18, output_MAC_73_19, 
		output_MAC_73_20, output_MAC_73_21, output_MAC_73_22, output_MAC_73_23, output_MAC_73_24, output_MAC_73_25, output_MAC_73_26, output_MAC_73_27, output_MAC_73_28, output_MAC_73_29, 
		output_MAC_73_30, output_MAC_73_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_74_0, output_MAC_74_1, output_MAC_74_2, output_MAC_74_3, output_MAC_74_4, output_MAC_74_5, output_MAC_74_6, output_MAC_74_7, output_MAC_74_8, output_MAC_74_9, 
		output_MAC_74_10, output_MAC_74_11, output_MAC_74_12, output_MAC_74_13, output_MAC_74_14, output_MAC_74_15, output_MAC_74_16, output_MAC_74_17, output_MAC_74_18, output_MAC_74_19, 
		output_MAC_74_20, output_MAC_74_21, output_MAC_74_22, output_MAC_74_23, output_MAC_74_24, output_MAC_74_25, output_MAC_74_26, output_MAC_74_27, output_MAC_74_28, output_MAC_74_29, 
		output_MAC_74_30, output_MAC_74_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_75_0, output_MAC_75_1, output_MAC_75_2, output_MAC_75_3, output_MAC_75_4, output_MAC_75_5, output_MAC_75_6, output_MAC_75_7, output_MAC_75_8, output_MAC_75_9, 
		output_MAC_75_10, output_MAC_75_11, output_MAC_75_12, output_MAC_75_13, output_MAC_75_14, output_MAC_75_15, output_MAC_75_16, output_MAC_75_17, output_MAC_75_18, output_MAC_75_19, 
		output_MAC_75_20, output_MAC_75_21, output_MAC_75_22, output_MAC_75_23, output_MAC_75_24, output_MAC_75_25, output_MAC_75_26, output_MAC_75_27, output_MAC_75_28, output_MAC_75_29, 
		output_MAC_75_30, output_MAC_75_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_76_0, output_MAC_76_1, output_MAC_76_2, output_MAC_76_3, output_MAC_76_4, output_MAC_76_5, output_MAC_76_6, output_MAC_76_7, output_MAC_76_8, output_MAC_76_9, 
		output_MAC_76_10, output_MAC_76_11, output_MAC_76_12, output_MAC_76_13, output_MAC_76_14, output_MAC_76_15, output_MAC_76_16, output_MAC_76_17, output_MAC_76_18, output_MAC_76_19, 
		output_MAC_76_20, output_MAC_76_21, output_MAC_76_22, output_MAC_76_23, output_MAC_76_24, output_MAC_76_25, output_MAC_76_26, output_MAC_76_27, output_MAC_76_28, output_MAC_76_29, 
		output_MAC_76_30, output_MAC_76_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_77_0, output_MAC_77_1, output_MAC_77_2, output_MAC_77_3, output_MAC_77_4, output_MAC_77_5, output_MAC_77_6, output_MAC_77_7, output_MAC_77_8, output_MAC_77_9, 
		output_MAC_77_10, output_MAC_77_11, output_MAC_77_12, output_MAC_77_13, output_MAC_77_14, output_MAC_77_15, output_MAC_77_16, output_MAC_77_17, output_MAC_77_18, output_MAC_77_19, 
		output_MAC_77_20, output_MAC_77_21, output_MAC_77_22, output_MAC_77_23, output_MAC_77_24, output_MAC_77_25, output_MAC_77_26, output_MAC_77_27, output_MAC_77_28, output_MAC_77_29, 
		output_MAC_77_30, output_MAC_77_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_78_0, output_MAC_78_1, output_MAC_78_2, output_MAC_78_3, output_MAC_78_4, output_MAC_78_5, output_MAC_78_6, output_MAC_78_7, output_MAC_78_8, output_MAC_78_9, 
		output_MAC_78_10, output_MAC_78_11, output_MAC_78_12, output_MAC_78_13, output_MAC_78_14, output_MAC_78_15, output_MAC_78_16, output_MAC_78_17, output_MAC_78_18, output_MAC_78_19, 
		output_MAC_78_20, output_MAC_78_21, output_MAC_78_22, output_MAC_78_23, output_MAC_78_24, output_MAC_78_25, output_MAC_78_26, output_MAC_78_27, output_MAC_78_28, output_MAC_78_29, 
		output_MAC_78_30, output_MAC_78_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_79_0, output_MAC_79_1, output_MAC_79_2, output_MAC_79_3, output_MAC_79_4, output_MAC_79_5, output_MAC_79_6, output_MAC_79_7, output_MAC_79_8, output_MAC_79_9, 
		output_MAC_79_10, output_MAC_79_11, output_MAC_79_12, output_MAC_79_13, output_MAC_79_14, output_MAC_79_15, output_MAC_79_16, output_MAC_79_17, output_MAC_79_18, output_MAC_79_19, 
		output_MAC_79_20, output_MAC_79_21, output_MAC_79_22, output_MAC_79_23, output_MAC_79_24, output_MAC_79_25, output_MAC_79_26, output_MAC_79_27, output_MAC_79_28, output_MAC_79_29, 
		output_MAC_79_30, output_MAC_79_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_80_0, output_MAC_80_1, output_MAC_80_2, output_MAC_80_3, output_MAC_80_4, output_MAC_80_5, output_MAC_80_6, output_MAC_80_7, output_MAC_80_8, output_MAC_80_9, 
		output_MAC_80_10, output_MAC_80_11, output_MAC_80_12, output_MAC_80_13, output_MAC_80_14, output_MAC_80_15, output_MAC_80_16, output_MAC_80_17, output_MAC_80_18, output_MAC_80_19, 
		output_MAC_80_20, output_MAC_80_21, output_MAC_80_22, output_MAC_80_23, output_MAC_80_24, output_MAC_80_25, output_MAC_80_26, output_MAC_80_27, output_MAC_80_28, output_MAC_80_29, 
		output_MAC_80_30, output_MAC_80_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_81_0, output_MAC_81_1, output_MAC_81_2, output_MAC_81_3, output_MAC_81_4, output_MAC_81_5, output_MAC_81_6, output_MAC_81_7, output_MAC_81_8, output_MAC_81_9, 
		output_MAC_81_10, output_MAC_81_11, output_MAC_81_12, output_MAC_81_13, output_MAC_81_14, output_MAC_81_15, output_MAC_81_16, output_MAC_81_17, output_MAC_81_18, output_MAC_81_19, 
		output_MAC_81_20, output_MAC_81_21, output_MAC_81_22, output_MAC_81_23, output_MAC_81_24, output_MAC_81_25, output_MAC_81_26, output_MAC_81_27, output_MAC_81_28, output_MAC_81_29, 
		output_MAC_81_30, output_MAC_81_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_82_0, output_MAC_82_1, output_MAC_82_2, output_MAC_82_3, output_MAC_82_4, output_MAC_82_5, output_MAC_82_6, output_MAC_82_7, output_MAC_82_8, output_MAC_82_9, 
		output_MAC_82_10, output_MAC_82_11, output_MAC_82_12, output_MAC_82_13, output_MAC_82_14, output_MAC_82_15, output_MAC_82_16, output_MAC_82_17, output_MAC_82_18, output_MAC_82_19, 
		output_MAC_82_20, output_MAC_82_21, output_MAC_82_22, output_MAC_82_23, output_MAC_82_24, output_MAC_82_25, output_MAC_82_26, output_MAC_82_27, output_MAC_82_28, output_MAC_82_29, 
		output_MAC_82_30, output_MAC_82_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_83_0, output_MAC_83_1, output_MAC_83_2, output_MAC_83_3, output_MAC_83_4, output_MAC_83_5, output_MAC_83_6, output_MAC_83_7, output_MAC_83_8, output_MAC_83_9, 
		output_MAC_83_10, output_MAC_83_11, output_MAC_83_12, output_MAC_83_13, output_MAC_83_14, output_MAC_83_15, output_MAC_83_16, output_MAC_83_17, output_MAC_83_18, output_MAC_83_19, 
		output_MAC_83_20, output_MAC_83_21, output_MAC_83_22, output_MAC_83_23, output_MAC_83_24, output_MAC_83_25, output_MAC_83_26, output_MAC_83_27, output_MAC_83_28, output_MAC_83_29, 
		output_MAC_83_30, output_MAC_83_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_84_0, output_MAC_84_1, output_MAC_84_2, output_MAC_84_3, output_MAC_84_4, output_MAC_84_5, output_MAC_84_6, output_MAC_84_7, output_MAC_84_8, output_MAC_84_9, 
		output_MAC_84_10, output_MAC_84_11, output_MAC_84_12, output_MAC_84_13, output_MAC_84_14, output_MAC_84_15, output_MAC_84_16, output_MAC_84_17, output_MAC_84_18, output_MAC_84_19, 
		output_MAC_84_20, output_MAC_84_21, output_MAC_84_22, output_MAC_84_23, output_MAC_84_24, output_MAC_84_25, output_MAC_84_26, output_MAC_84_27, output_MAC_84_28, output_MAC_84_29, 
		output_MAC_84_30, output_MAC_84_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_85_0, output_MAC_85_1, output_MAC_85_2, output_MAC_85_3, output_MAC_85_4, output_MAC_85_5, output_MAC_85_6, output_MAC_85_7, output_MAC_85_8, output_MAC_85_9, 
		output_MAC_85_10, output_MAC_85_11, output_MAC_85_12, output_MAC_85_13, output_MAC_85_14, output_MAC_85_15, output_MAC_85_16, output_MAC_85_17, output_MAC_85_18, output_MAC_85_19, 
		output_MAC_85_20, output_MAC_85_21, output_MAC_85_22, output_MAC_85_23, output_MAC_85_24, output_MAC_85_25, output_MAC_85_26, output_MAC_85_27, output_MAC_85_28, output_MAC_85_29, 
		output_MAC_85_30, output_MAC_85_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_86_0, output_MAC_86_1, output_MAC_86_2, output_MAC_86_3, output_MAC_86_4, output_MAC_86_5, output_MAC_86_6, output_MAC_86_7, output_MAC_86_8, output_MAC_86_9, 
		output_MAC_86_10, output_MAC_86_11, output_MAC_86_12, output_MAC_86_13, output_MAC_86_14, output_MAC_86_15, output_MAC_86_16, output_MAC_86_17, output_MAC_86_18, output_MAC_86_19, 
		output_MAC_86_20, output_MAC_86_21, output_MAC_86_22, output_MAC_86_23, output_MAC_86_24, output_MAC_86_25, output_MAC_86_26, output_MAC_86_27, output_MAC_86_28, output_MAC_86_29, 
		output_MAC_86_30, output_MAC_86_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_87_0, output_MAC_87_1, output_MAC_87_2, output_MAC_87_3, output_MAC_87_4, output_MAC_87_5, output_MAC_87_6, output_MAC_87_7, output_MAC_87_8, output_MAC_87_9, 
		output_MAC_87_10, output_MAC_87_11, output_MAC_87_12, output_MAC_87_13, output_MAC_87_14, output_MAC_87_15, output_MAC_87_16, output_MAC_87_17, output_MAC_87_18, output_MAC_87_19, 
		output_MAC_87_20, output_MAC_87_21, output_MAC_87_22, output_MAC_87_23, output_MAC_87_24, output_MAC_87_25, output_MAC_87_26, output_MAC_87_27, output_MAC_87_28, output_MAC_87_29, 
		output_MAC_87_30, output_MAC_87_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_88_0, output_MAC_88_1, output_MAC_88_2, output_MAC_88_3, output_MAC_88_4, output_MAC_88_5, output_MAC_88_6, output_MAC_88_7, output_MAC_88_8, output_MAC_88_9, 
		output_MAC_88_10, output_MAC_88_11, output_MAC_88_12, output_MAC_88_13, output_MAC_88_14, output_MAC_88_15, output_MAC_88_16, output_MAC_88_17, output_MAC_88_18, output_MAC_88_19, 
		output_MAC_88_20, output_MAC_88_21, output_MAC_88_22, output_MAC_88_23, output_MAC_88_24, output_MAC_88_25, output_MAC_88_26, output_MAC_88_27, output_MAC_88_28, output_MAC_88_29, 
		output_MAC_88_30, output_MAC_88_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_89_0, output_MAC_89_1, output_MAC_89_2, output_MAC_89_3, output_MAC_89_4, output_MAC_89_5, output_MAC_89_6, output_MAC_89_7, output_MAC_89_8, output_MAC_89_9, 
		output_MAC_89_10, output_MAC_89_11, output_MAC_89_12, output_MAC_89_13, output_MAC_89_14, output_MAC_89_15, output_MAC_89_16, output_MAC_89_17, output_MAC_89_18, output_MAC_89_19, 
		output_MAC_89_20, output_MAC_89_21, output_MAC_89_22, output_MAC_89_23, output_MAC_89_24, output_MAC_89_25, output_MAC_89_26, output_MAC_89_27, output_MAC_89_28, output_MAC_89_29, 
		output_MAC_89_30, output_MAC_89_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_90_0, output_MAC_90_1, output_MAC_90_2, output_MAC_90_3, output_MAC_90_4, output_MAC_90_5, output_MAC_90_6, output_MAC_90_7, output_MAC_90_8, output_MAC_90_9, 
		output_MAC_90_10, output_MAC_90_11, output_MAC_90_12, output_MAC_90_13, output_MAC_90_14, output_MAC_90_15, output_MAC_90_16, output_MAC_90_17, output_MAC_90_18, output_MAC_90_19, 
		output_MAC_90_20, output_MAC_90_21, output_MAC_90_22, output_MAC_90_23, output_MAC_90_24, output_MAC_90_25, output_MAC_90_26, output_MAC_90_27, output_MAC_90_28, output_MAC_90_29, 
		output_MAC_90_30, output_MAC_90_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_91_0, output_MAC_91_1, output_MAC_91_2, output_MAC_91_3, output_MAC_91_4, output_MAC_91_5, output_MAC_91_6, output_MAC_91_7, output_MAC_91_8, output_MAC_91_9, 
		output_MAC_91_10, output_MAC_91_11, output_MAC_91_12, output_MAC_91_13, output_MAC_91_14, output_MAC_91_15, output_MAC_91_16, output_MAC_91_17, output_MAC_91_18, output_MAC_91_19, 
		output_MAC_91_20, output_MAC_91_21, output_MAC_91_22, output_MAC_91_23, output_MAC_91_24, output_MAC_91_25, output_MAC_91_26, output_MAC_91_27, output_MAC_91_28, output_MAC_91_29, 
		output_MAC_91_30, output_MAC_91_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_92_0, output_MAC_92_1, output_MAC_92_2, output_MAC_92_3, output_MAC_92_4, output_MAC_92_5, output_MAC_92_6, output_MAC_92_7, output_MAC_92_8, output_MAC_92_9, 
		output_MAC_92_10, output_MAC_92_11, output_MAC_92_12, output_MAC_92_13, output_MAC_92_14, output_MAC_92_15, output_MAC_92_16, output_MAC_92_17, output_MAC_92_18, output_MAC_92_19, 
		output_MAC_92_20, output_MAC_92_21, output_MAC_92_22, output_MAC_92_23, output_MAC_92_24, output_MAC_92_25, output_MAC_92_26, output_MAC_92_27, output_MAC_92_28, output_MAC_92_29, 
		output_MAC_92_30, output_MAC_92_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_93_0, output_MAC_93_1, output_MAC_93_2, output_MAC_93_3, output_MAC_93_4, output_MAC_93_5, output_MAC_93_6, output_MAC_93_7, output_MAC_93_8, output_MAC_93_9, 
		output_MAC_93_10, output_MAC_93_11, output_MAC_93_12, output_MAC_93_13, output_MAC_93_14, output_MAC_93_15, output_MAC_93_16, output_MAC_93_17, output_MAC_93_18, output_MAC_93_19, 
		output_MAC_93_20, output_MAC_93_21, output_MAC_93_22, output_MAC_93_23, output_MAC_93_24, output_MAC_93_25, output_MAC_93_26, output_MAC_93_27, output_MAC_93_28, output_MAC_93_29, 
		output_MAC_93_30, output_MAC_93_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_94_0, output_MAC_94_1, output_MAC_94_2, output_MAC_94_3, output_MAC_94_4, output_MAC_94_5, output_MAC_94_6, output_MAC_94_7, output_MAC_94_8, output_MAC_94_9, 
		output_MAC_94_10, output_MAC_94_11, output_MAC_94_12, output_MAC_94_13, output_MAC_94_14, output_MAC_94_15, output_MAC_94_16, output_MAC_94_17, output_MAC_94_18, output_MAC_94_19, 
		output_MAC_94_20, output_MAC_94_21, output_MAC_94_22, output_MAC_94_23, output_MAC_94_24, output_MAC_94_25, output_MAC_94_26, output_MAC_94_27, output_MAC_94_28, output_MAC_94_29, 
		output_MAC_94_30, output_MAC_94_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_95_0, output_MAC_95_1, output_MAC_95_2, output_MAC_95_3, output_MAC_95_4, output_MAC_95_5, output_MAC_95_6, output_MAC_95_7, output_MAC_95_8, output_MAC_95_9, 
		output_MAC_95_10, output_MAC_95_11, output_MAC_95_12, output_MAC_95_13, output_MAC_95_14, output_MAC_95_15, output_MAC_95_16, output_MAC_95_17, output_MAC_95_18, output_MAC_95_19, 
		output_MAC_95_20, output_MAC_95_21, output_MAC_95_22, output_MAC_95_23, output_MAC_95_24, output_MAC_95_25, output_MAC_95_26, output_MAC_95_27, output_MAC_95_28, output_MAC_95_29, 
		output_MAC_95_30, output_MAC_95_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_96_0, output_MAC_96_1, output_MAC_96_2, output_MAC_96_3, output_MAC_96_4, output_MAC_96_5, output_MAC_96_6, output_MAC_96_7, output_MAC_96_8, output_MAC_96_9, 
		output_MAC_96_10, output_MAC_96_11, output_MAC_96_12, output_MAC_96_13, output_MAC_96_14, output_MAC_96_15, output_MAC_96_16, output_MAC_96_17, output_MAC_96_18, output_MAC_96_19, 
		output_MAC_96_20, output_MAC_96_21, output_MAC_96_22, output_MAC_96_23, output_MAC_96_24, output_MAC_96_25, output_MAC_96_26, output_MAC_96_27, output_MAC_96_28, output_MAC_96_29, 
		output_MAC_96_30, output_MAC_96_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_97_0, output_MAC_97_1, output_MAC_97_2, output_MAC_97_3, output_MAC_97_4, output_MAC_97_5, output_MAC_97_6, output_MAC_97_7, output_MAC_97_8, output_MAC_97_9, 
		output_MAC_97_10, output_MAC_97_11, output_MAC_97_12, output_MAC_97_13, output_MAC_97_14, output_MAC_97_15, output_MAC_97_16, output_MAC_97_17, output_MAC_97_18, output_MAC_97_19, 
		output_MAC_97_20, output_MAC_97_21, output_MAC_97_22, output_MAC_97_23, output_MAC_97_24, output_MAC_97_25, output_MAC_97_26, output_MAC_97_27, output_MAC_97_28, output_MAC_97_29, 
		output_MAC_97_30, output_MAC_97_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_98_0, output_MAC_98_1, output_MAC_98_2, output_MAC_98_3, output_MAC_98_4, output_MAC_98_5, output_MAC_98_6, output_MAC_98_7, output_MAC_98_8, output_MAC_98_9, 
		output_MAC_98_10, output_MAC_98_11, output_MAC_98_12, output_MAC_98_13, output_MAC_98_14, output_MAC_98_15, output_MAC_98_16, output_MAC_98_17, output_MAC_98_18, output_MAC_98_19, 
		output_MAC_98_20, output_MAC_98_21, output_MAC_98_22, output_MAC_98_23, output_MAC_98_24, output_MAC_98_25, output_MAC_98_26, output_MAC_98_27, output_MAC_98_28, output_MAC_98_29, 
		output_MAC_98_30, output_MAC_98_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_99_0, output_MAC_99_1, output_MAC_99_2, output_MAC_99_3, output_MAC_99_4, output_MAC_99_5, output_MAC_99_6, output_MAC_99_7, output_MAC_99_8, output_MAC_99_9, 
		output_MAC_99_10, output_MAC_99_11, output_MAC_99_12, output_MAC_99_13, output_MAC_99_14, output_MAC_99_15, output_MAC_99_16, output_MAC_99_17, output_MAC_99_18, output_MAC_99_19, 
		output_MAC_99_20, output_MAC_99_21, output_MAC_99_22, output_MAC_99_23, output_MAC_99_24, output_MAC_99_25, output_MAC_99_26, output_MAC_99_27, output_MAC_99_28, output_MAC_99_29, 
		output_MAC_99_30, output_MAC_99_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_100_0, output_MAC_100_1, output_MAC_100_2, output_MAC_100_3, output_MAC_100_4, output_MAC_100_5, output_MAC_100_6, output_MAC_100_7, output_MAC_100_8, output_MAC_100_9, 
		output_MAC_100_10, output_MAC_100_11, output_MAC_100_12, output_MAC_100_13, output_MAC_100_14, output_MAC_100_15, output_MAC_100_16, output_MAC_100_17, output_MAC_100_18, output_MAC_100_19, 
		output_MAC_100_20, output_MAC_100_21, output_MAC_100_22, output_MAC_100_23, output_MAC_100_24, output_MAC_100_25, output_MAC_100_26, output_MAC_100_27, output_MAC_100_28, output_MAC_100_29, 
		output_MAC_100_30, output_MAC_100_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_101_0, output_MAC_101_1, output_MAC_101_2, output_MAC_101_3, output_MAC_101_4, output_MAC_101_5, output_MAC_101_6, output_MAC_101_7, output_MAC_101_8, output_MAC_101_9, 
		output_MAC_101_10, output_MAC_101_11, output_MAC_101_12, output_MAC_101_13, output_MAC_101_14, output_MAC_101_15, output_MAC_101_16, output_MAC_101_17, output_MAC_101_18, output_MAC_101_19, 
		output_MAC_101_20, output_MAC_101_21, output_MAC_101_22, output_MAC_101_23, output_MAC_101_24, output_MAC_101_25, output_MAC_101_26, output_MAC_101_27, output_MAC_101_28, output_MAC_101_29, 
		output_MAC_101_30, output_MAC_101_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_102_0, output_MAC_102_1, output_MAC_102_2, output_MAC_102_3, output_MAC_102_4, output_MAC_102_5, output_MAC_102_6, output_MAC_102_7, output_MAC_102_8, output_MAC_102_9, 
		output_MAC_102_10, output_MAC_102_11, output_MAC_102_12, output_MAC_102_13, output_MAC_102_14, output_MAC_102_15, output_MAC_102_16, output_MAC_102_17, output_MAC_102_18, output_MAC_102_19, 
		output_MAC_102_20, output_MAC_102_21, output_MAC_102_22, output_MAC_102_23, output_MAC_102_24, output_MAC_102_25, output_MAC_102_26, output_MAC_102_27, output_MAC_102_28, output_MAC_102_29, 
		output_MAC_102_30, output_MAC_102_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_103_0, output_MAC_103_1, output_MAC_103_2, output_MAC_103_3, output_MAC_103_4, output_MAC_103_5, output_MAC_103_6, output_MAC_103_7, output_MAC_103_8, output_MAC_103_9, 
		output_MAC_103_10, output_MAC_103_11, output_MAC_103_12, output_MAC_103_13, output_MAC_103_14, output_MAC_103_15, output_MAC_103_16, output_MAC_103_17, output_MAC_103_18, output_MAC_103_19, 
		output_MAC_103_20, output_MAC_103_21, output_MAC_103_22, output_MAC_103_23, output_MAC_103_24, output_MAC_103_25, output_MAC_103_26, output_MAC_103_27, output_MAC_103_28, output_MAC_103_29, 
		output_MAC_103_30, output_MAC_103_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_104_0, output_MAC_104_1, output_MAC_104_2, output_MAC_104_3, output_MAC_104_4, output_MAC_104_5, output_MAC_104_6, output_MAC_104_7, output_MAC_104_8, output_MAC_104_9, 
		output_MAC_104_10, output_MAC_104_11, output_MAC_104_12, output_MAC_104_13, output_MAC_104_14, output_MAC_104_15, output_MAC_104_16, output_MAC_104_17, output_MAC_104_18, output_MAC_104_19, 
		output_MAC_104_20, output_MAC_104_21, output_MAC_104_22, output_MAC_104_23, output_MAC_104_24, output_MAC_104_25, output_MAC_104_26, output_MAC_104_27, output_MAC_104_28, output_MAC_104_29, 
		output_MAC_104_30, output_MAC_104_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_105_0, output_MAC_105_1, output_MAC_105_2, output_MAC_105_3, output_MAC_105_4, output_MAC_105_5, output_MAC_105_6, output_MAC_105_7, output_MAC_105_8, output_MAC_105_9, 
		output_MAC_105_10, output_MAC_105_11, output_MAC_105_12, output_MAC_105_13, output_MAC_105_14, output_MAC_105_15, output_MAC_105_16, output_MAC_105_17, output_MAC_105_18, output_MAC_105_19, 
		output_MAC_105_20, output_MAC_105_21, output_MAC_105_22, output_MAC_105_23, output_MAC_105_24, output_MAC_105_25, output_MAC_105_26, output_MAC_105_27, output_MAC_105_28, output_MAC_105_29, 
		output_MAC_105_30, output_MAC_105_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_106_0, output_MAC_106_1, output_MAC_106_2, output_MAC_106_3, output_MAC_106_4, output_MAC_106_5, output_MAC_106_6, output_MAC_106_7, output_MAC_106_8, output_MAC_106_9, 
		output_MAC_106_10, output_MAC_106_11, output_MAC_106_12, output_MAC_106_13, output_MAC_106_14, output_MAC_106_15, output_MAC_106_16, output_MAC_106_17, output_MAC_106_18, output_MAC_106_19, 
		output_MAC_106_20, output_MAC_106_21, output_MAC_106_22, output_MAC_106_23, output_MAC_106_24, output_MAC_106_25, output_MAC_106_26, output_MAC_106_27, output_MAC_106_28, output_MAC_106_29, 
		output_MAC_106_30, output_MAC_106_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_107_0, output_MAC_107_1, output_MAC_107_2, output_MAC_107_3, output_MAC_107_4, output_MAC_107_5, output_MAC_107_6, output_MAC_107_7, output_MAC_107_8, output_MAC_107_9, 
		output_MAC_107_10, output_MAC_107_11, output_MAC_107_12, output_MAC_107_13, output_MAC_107_14, output_MAC_107_15, output_MAC_107_16, output_MAC_107_17, output_MAC_107_18, output_MAC_107_19, 
		output_MAC_107_20, output_MAC_107_21, output_MAC_107_22, output_MAC_107_23, output_MAC_107_24, output_MAC_107_25, output_MAC_107_26, output_MAC_107_27, output_MAC_107_28, output_MAC_107_29, 
		output_MAC_107_30, output_MAC_107_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_108_0, output_MAC_108_1, output_MAC_108_2, output_MAC_108_3, output_MAC_108_4, output_MAC_108_5, output_MAC_108_6, output_MAC_108_7, output_MAC_108_8, output_MAC_108_9, 
		output_MAC_108_10, output_MAC_108_11, output_MAC_108_12, output_MAC_108_13, output_MAC_108_14, output_MAC_108_15, output_MAC_108_16, output_MAC_108_17, output_MAC_108_18, output_MAC_108_19, 
		output_MAC_108_20, output_MAC_108_21, output_MAC_108_22, output_MAC_108_23, output_MAC_108_24, output_MAC_108_25, output_MAC_108_26, output_MAC_108_27, output_MAC_108_28, output_MAC_108_29, 
		output_MAC_108_30, output_MAC_108_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_109_0, output_MAC_109_1, output_MAC_109_2, output_MAC_109_3, output_MAC_109_4, output_MAC_109_5, output_MAC_109_6, output_MAC_109_7, output_MAC_109_8, output_MAC_109_9, 
		output_MAC_109_10, output_MAC_109_11, output_MAC_109_12, output_MAC_109_13, output_MAC_109_14, output_MAC_109_15, output_MAC_109_16, output_MAC_109_17, output_MAC_109_18, output_MAC_109_19, 
		output_MAC_109_20, output_MAC_109_21, output_MAC_109_22, output_MAC_109_23, output_MAC_109_24, output_MAC_109_25, output_MAC_109_26, output_MAC_109_27, output_MAC_109_28, output_MAC_109_29, 
		output_MAC_109_30, output_MAC_109_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_110_0, output_MAC_110_1, output_MAC_110_2, output_MAC_110_3, output_MAC_110_4, output_MAC_110_5, output_MAC_110_6, output_MAC_110_7, output_MAC_110_8, output_MAC_110_9, 
		output_MAC_110_10, output_MAC_110_11, output_MAC_110_12, output_MAC_110_13, output_MAC_110_14, output_MAC_110_15, output_MAC_110_16, output_MAC_110_17, output_MAC_110_18, output_MAC_110_19, 
		output_MAC_110_20, output_MAC_110_21, output_MAC_110_22, output_MAC_110_23, output_MAC_110_24, output_MAC_110_25, output_MAC_110_26, output_MAC_110_27, output_MAC_110_28, output_MAC_110_29, 
		output_MAC_110_30, output_MAC_110_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_111_0, output_MAC_111_1, output_MAC_111_2, output_MAC_111_3, output_MAC_111_4, output_MAC_111_5, output_MAC_111_6, output_MAC_111_7, output_MAC_111_8, output_MAC_111_9, 
		output_MAC_111_10, output_MAC_111_11, output_MAC_111_12, output_MAC_111_13, output_MAC_111_14, output_MAC_111_15, output_MAC_111_16, output_MAC_111_17, output_MAC_111_18, output_MAC_111_19, 
		output_MAC_111_20, output_MAC_111_21, output_MAC_111_22, output_MAC_111_23, output_MAC_111_24, output_MAC_111_25, output_MAC_111_26, output_MAC_111_27, output_MAC_111_28, output_MAC_111_29, 
		output_MAC_111_30, output_MAC_111_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_112_0, output_MAC_112_1, output_MAC_112_2, output_MAC_112_3, output_MAC_112_4, output_MAC_112_5, output_MAC_112_6, output_MAC_112_7, output_MAC_112_8, output_MAC_112_9, 
		output_MAC_112_10, output_MAC_112_11, output_MAC_112_12, output_MAC_112_13, output_MAC_112_14, output_MAC_112_15, output_MAC_112_16, output_MAC_112_17, output_MAC_112_18, output_MAC_112_19, 
		output_MAC_112_20, output_MAC_112_21, output_MAC_112_22, output_MAC_112_23, output_MAC_112_24, output_MAC_112_25, output_MAC_112_26, output_MAC_112_27, output_MAC_112_28, output_MAC_112_29, 
		output_MAC_112_30, output_MAC_112_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_113_0, output_MAC_113_1, output_MAC_113_2, output_MAC_113_3, output_MAC_113_4, output_MAC_113_5, output_MAC_113_6, output_MAC_113_7, output_MAC_113_8, output_MAC_113_9, 
		output_MAC_113_10, output_MAC_113_11, output_MAC_113_12, output_MAC_113_13, output_MAC_113_14, output_MAC_113_15, output_MAC_113_16, output_MAC_113_17, output_MAC_113_18, output_MAC_113_19, 
		output_MAC_113_20, output_MAC_113_21, output_MAC_113_22, output_MAC_113_23, output_MAC_113_24, output_MAC_113_25, output_MAC_113_26, output_MAC_113_27, output_MAC_113_28, output_MAC_113_29, 
		output_MAC_113_30, output_MAC_113_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_114_0, output_MAC_114_1, output_MAC_114_2, output_MAC_114_3, output_MAC_114_4, output_MAC_114_5, output_MAC_114_6, output_MAC_114_7, output_MAC_114_8, output_MAC_114_9, 
		output_MAC_114_10, output_MAC_114_11, output_MAC_114_12, output_MAC_114_13, output_MAC_114_14, output_MAC_114_15, output_MAC_114_16, output_MAC_114_17, output_MAC_114_18, output_MAC_114_19, 
		output_MAC_114_20, output_MAC_114_21, output_MAC_114_22, output_MAC_114_23, output_MAC_114_24, output_MAC_114_25, output_MAC_114_26, output_MAC_114_27, output_MAC_114_28, output_MAC_114_29, 
		output_MAC_114_30, output_MAC_114_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_115_0, output_MAC_115_1, output_MAC_115_2, output_MAC_115_3, output_MAC_115_4, output_MAC_115_5, output_MAC_115_6, output_MAC_115_7, output_MAC_115_8, output_MAC_115_9, 
		output_MAC_115_10, output_MAC_115_11, output_MAC_115_12, output_MAC_115_13, output_MAC_115_14, output_MAC_115_15, output_MAC_115_16, output_MAC_115_17, output_MAC_115_18, output_MAC_115_19, 
		output_MAC_115_20, output_MAC_115_21, output_MAC_115_22, output_MAC_115_23, output_MAC_115_24, output_MAC_115_25, output_MAC_115_26, output_MAC_115_27, output_MAC_115_28, output_MAC_115_29, 
		output_MAC_115_30, output_MAC_115_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_116_0, output_MAC_116_1, output_MAC_116_2, output_MAC_116_3, output_MAC_116_4, output_MAC_116_5, output_MAC_116_6, output_MAC_116_7, output_MAC_116_8, output_MAC_116_9, 
		output_MAC_116_10, output_MAC_116_11, output_MAC_116_12, output_MAC_116_13, output_MAC_116_14, output_MAC_116_15, output_MAC_116_16, output_MAC_116_17, output_MAC_116_18, output_MAC_116_19, 
		output_MAC_116_20, output_MAC_116_21, output_MAC_116_22, output_MAC_116_23, output_MAC_116_24, output_MAC_116_25, output_MAC_116_26, output_MAC_116_27, output_MAC_116_28, output_MAC_116_29, 
		output_MAC_116_30, output_MAC_116_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_117_0, output_MAC_117_1, output_MAC_117_2, output_MAC_117_3, output_MAC_117_4, output_MAC_117_5, output_MAC_117_6, output_MAC_117_7, output_MAC_117_8, output_MAC_117_9, 
		output_MAC_117_10, output_MAC_117_11, output_MAC_117_12, output_MAC_117_13, output_MAC_117_14, output_MAC_117_15, output_MAC_117_16, output_MAC_117_17, output_MAC_117_18, output_MAC_117_19, 
		output_MAC_117_20, output_MAC_117_21, output_MAC_117_22, output_MAC_117_23, output_MAC_117_24, output_MAC_117_25, output_MAC_117_26, output_MAC_117_27, output_MAC_117_28, output_MAC_117_29, 
		output_MAC_117_30, output_MAC_117_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_118_0, output_MAC_118_1, output_MAC_118_2, output_MAC_118_3, output_MAC_118_4, output_MAC_118_5, output_MAC_118_6, output_MAC_118_7, output_MAC_118_8, output_MAC_118_9, 
		output_MAC_118_10, output_MAC_118_11, output_MAC_118_12, output_MAC_118_13, output_MAC_118_14, output_MAC_118_15, output_MAC_118_16, output_MAC_118_17, output_MAC_118_18, output_MAC_118_19, 
		output_MAC_118_20, output_MAC_118_21, output_MAC_118_22, output_MAC_118_23, output_MAC_118_24, output_MAC_118_25, output_MAC_118_26, output_MAC_118_27, output_MAC_118_28, output_MAC_118_29, 
		output_MAC_118_30, output_MAC_118_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_119_0, output_MAC_119_1, output_MAC_119_2, output_MAC_119_3, output_MAC_119_4, output_MAC_119_5, output_MAC_119_6, output_MAC_119_7, output_MAC_119_8, output_MAC_119_9, 
		output_MAC_119_10, output_MAC_119_11, output_MAC_119_12, output_MAC_119_13, output_MAC_119_14, output_MAC_119_15, output_MAC_119_16, output_MAC_119_17, output_MAC_119_18, output_MAC_119_19, 
		output_MAC_119_20, output_MAC_119_21, output_MAC_119_22, output_MAC_119_23, output_MAC_119_24, output_MAC_119_25, output_MAC_119_26, output_MAC_119_27, output_MAC_119_28, output_MAC_119_29, 
		output_MAC_119_30, output_MAC_119_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_120_0, output_MAC_120_1, output_MAC_120_2, output_MAC_120_3, output_MAC_120_4, output_MAC_120_5, output_MAC_120_6, output_MAC_120_7, output_MAC_120_8, output_MAC_120_9, 
		output_MAC_120_10, output_MAC_120_11, output_MAC_120_12, output_MAC_120_13, output_MAC_120_14, output_MAC_120_15, output_MAC_120_16, output_MAC_120_17, output_MAC_120_18, output_MAC_120_19, 
		output_MAC_120_20, output_MAC_120_21, output_MAC_120_22, output_MAC_120_23, output_MAC_120_24, output_MAC_120_25, output_MAC_120_26, output_MAC_120_27, output_MAC_120_28, output_MAC_120_29, 
		output_MAC_120_30, output_MAC_120_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_121_0, output_MAC_121_1, output_MAC_121_2, output_MAC_121_3, output_MAC_121_4, output_MAC_121_5, output_MAC_121_6, output_MAC_121_7, output_MAC_121_8, output_MAC_121_9, 
		output_MAC_121_10, output_MAC_121_11, output_MAC_121_12, output_MAC_121_13, output_MAC_121_14, output_MAC_121_15, output_MAC_121_16, output_MAC_121_17, output_MAC_121_18, output_MAC_121_19, 
		output_MAC_121_20, output_MAC_121_21, output_MAC_121_22, output_MAC_121_23, output_MAC_121_24, output_MAC_121_25, output_MAC_121_26, output_MAC_121_27, output_MAC_121_28, output_MAC_121_29, 
		output_MAC_121_30, output_MAC_121_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_122_0, output_MAC_122_1, output_MAC_122_2, output_MAC_122_3, output_MAC_122_4, output_MAC_122_5, output_MAC_122_6, output_MAC_122_7, output_MAC_122_8, output_MAC_122_9, 
		output_MAC_122_10, output_MAC_122_11, output_MAC_122_12, output_MAC_122_13, output_MAC_122_14, output_MAC_122_15, output_MAC_122_16, output_MAC_122_17, output_MAC_122_18, output_MAC_122_19, 
		output_MAC_122_20, output_MAC_122_21, output_MAC_122_22, output_MAC_122_23, output_MAC_122_24, output_MAC_122_25, output_MAC_122_26, output_MAC_122_27, output_MAC_122_28, output_MAC_122_29, 
		output_MAC_122_30, output_MAC_122_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_123_0, output_MAC_123_1, output_MAC_123_2, output_MAC_123_3, output_MAC_123_4, output_MAC_123_5, output_MAC_123_6, output_MAC_123_7, output_MAC_123_8, output_MAC_123_9, 
		output_MAC_123_10, output_MAC_123_11, output_MAC_123_12, output_MAC_123_13, output_MAC_123_14, output_MAC_123_15, output_MAC_123_16, output_MAC_123_17, output_MAC_123_18, output_MAC_123_19, 
		output_MAC_123_20, output_MAC_123_21, output_MAC_123_22, output_MAC_123_23, output_MAC_123_24, output_MAC_123_25, output_MAC_123_26, output_MAC_123_27, output_MAC_123_28, output_MAC_123_29, 
		output_MAC_123_30, output_MAC_123_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_124_0, output_MAC_124_1, output_MAC_124_2, output_MAC_124_3, output_MAC_124_4, output_MAC_124_5, output_MAC_124_6, output_MAC_124_7, output_MAC_124_8, output_MAC_124_9, 
		output_MAC_124_10, output_MAC_124_11, output_MAC_124_12, output_MAC_124_13, output_MAC_124_14, output_MAC_124_15, output_MAC_124_16, output_MAC_124_17, output_MAC_124_18, output_MAC_124_19, 
		output_MAC_124_20, output_MAC_124_21, output_MAC_124_22, output_MAC_124_23, output_MAC_124_24, output_MAC_124_25, output_MAC_124_26, output_MAC_124_27, output_MAC_124_28, output_MAC_124_29, 
		output_MAC_124_30, output_MAC_124_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_125_0, output_MAC_125_1, output_MAC_125_2, output_MAC_125_3, output_MAC_125_4, output_MAC_125_5, output_MAC_125_6, output_MAC_125_7, output_MAC_125_8, output_MAC_125_9, 
		output_MAC_125_10, output_MAC_125_11, output_MAC_125_12, output_MAC_125_13, output_MAC_125_14, output_MAC_125_15, output_MAC_125_16, output_MAC_125_17, output_MAC_125_18, output_MAC_125_19, 
		output_MAC_125_20, output_MAC_125_21, output_MAC_125_22, output_MAC_125_23, output_MAC_125_24, output_MAC_125_25, output_MAC_125_26, output_MAC_125_27, output_MAC_125_28, output_MAC_125_29, 
		output_MAC_125_30, output_MAC_125_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_126_0, output_MAC_126_1, output_MAC_126_2, output_MAC_126_3, output_MAC_126_4, output_MAC_126_5, output_MAC_126_6, output_MAC_126_7, output_MAC_126_8, output_MAC_126_9, 
		output_MAC_126_10, output_MAC_126_11, output_MAC_126_12, output_MAC_126_13, output_MAC_126_14, output_MAC_126_15, output_MAC_126_16, output_MAC_126_17, output_MAC_126_18, output_MAC_126_19, 
		output_MAC_126_20, output_MAC_126_21, output_MAC_126_22, output_MAC_126_23, output_MAC_126_24, output_MAC_126_25, output_MAC_126_26, output_MAC_126_27, output_MAC_126_28, output_MAC_126_29, 
		output_MAC_126_30, output_MAC_126_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_127_0, output_MAC_127_1, output_MAC_127_2, output_MAC_127_3, output_MAC_127_4, output_MAC_127_5, output_MAC_127_6, output_MAC_127_7, output_MAC_127_8, output_MAC_127_9, 
		output_MAC_127_10, output_MAC_127_11, output_MAC_127_12, output_MAC_127_13, output_MAC_127_14, output_MAC_127_15, output_MAC_127_16, output_MAC_127_17, output_MAC_127_18, output_MAC_127_19, 
		output_MAC_127_20, output_MAC_127_21, output_MAC_127_22, output_MAC_127_23, output_MAC_127_24, output_MAC_127_25, output_MAC_127_26, output_MAC_127_27, output_MAC_127_28, output_MAC_127_29, 
		output_MAC_127_30, output_MAC_127_31: STD_LOGIC_VECTOR(31 downto 0);

BEGIN

	input_row_0_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_0, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_0);
	input_row_1_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_1, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_1);
	input_row_2_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_2, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_2);
	input_row_3_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_3, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_3);
	input_row_4_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_4, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_4);
	input_row_5_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_5, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_5);
	input_row_6_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_6, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_6);
	input_row_7_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_7, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_7);
	input_row_8_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_8, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_8);
	input_row_9_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_9, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_9);
	input_row_10_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_10, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_10);
	input_row_11_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_11, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_11);
	input_row_12_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_12, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_12);
	input_row_13_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_13, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_13);
	input_row_14_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_14, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_14);
	input_row_15_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_15, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_15);
	input_row_16_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_16, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_16);
	input_row_17_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_17, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_17);
	input_row_18_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_18, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_18);
	input_row_19_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_19, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_19);
	input_row_20_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_20, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_20);
	input_row_21_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_21, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_21);
	input_row_22_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_22, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_22);
	input_row_23_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_23, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_23);
	input_row_24_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_24, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_24);
	input_row_25_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_25, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_25);
	input_row_26_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_26, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_26);
	input_row_27_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_27, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_27);
	input_row_28_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_28, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_28);
	input_row_29_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_29, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_29);
	input_row_30_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_30, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_30);
	input_row_31_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_31, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_31);
	input_row_32_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_32, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_32);
	input_row_33_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_33, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_33);
	input_row_34_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_34, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_34);
	input_row_35_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_35, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_35);
	input_row_36_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_36, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_36);
	input_row_37_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_37, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_37);
	input_row_38_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_38, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_38);
	input_row_39_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_39, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_39);
	input_row_40_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_40, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_40);
	input_row_41_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_41, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_41);
	input_row_42_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_42, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_42);
	input_row_43_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_43, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_43);
	input_row_44_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_44, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_44);
	input_row_45_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_45, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_45);
	input_row_46_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_46, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_46);
	input_row_47_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_47, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_47);
	input_row_48_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_48, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_48);
	input_row_49_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_49, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_49);
	input_row_50_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_50, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_50);
	input_row_51_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_51, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_51);
	input_row_52_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_52, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_52);
	input_row_53_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_53, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_53);
	input_row_54_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_54, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_54);
	input_row_55_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_55, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_55);
	input_row_56_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_56, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_56);
	input_row_57_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_57, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_57);
	input_row_58_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_58, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_58);
	input_row_59_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_59, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_59);
	input_row_60_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_60, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_60);
	input_row_61_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_61, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_61);
	input_row_62_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_62, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_62);
	input_row_63_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_63, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_63);
	input_row_64_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_64, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_64);
	input_row_65_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_65, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_65);
	input_row_66_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_66, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_66);
	input_row_67_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_67, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_67);
	input_row_68_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_68, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_68);
	input_row_69_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_69, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_69);
	input_row_70_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_70, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_70);
	input_row_71_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_71, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_71);
	input_row_72_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_72, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_72);
	input_row_73_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_73, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_73);
	input_row_74_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_74, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_74);
	input_row_75_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_75, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_75);
	input_row_76_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_76, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_76);
	input_row_77_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_77, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_77);
	input_row_78_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_78, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_78);
	input_row_79_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_79, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_79);
	input_row_80_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_80, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_80);
	input_row_81_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_81, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_81);
	input_row_82_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_82, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_82);
	input_row_83_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_83, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_83);
	input_row_84_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_84, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_84);
	input_row_85_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_85, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_85);
	input_row_86_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_86, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_86);
	input_row_87_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_87, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_87);
	input_row_88_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_88, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_88);
	input_row_89_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_89, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_89);
	input_row_90_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_90, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_90);
	input_row_91_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_91, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_91);
	input_row_92_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_92, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_92);
	input_row_93_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_93, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_93);
	input_row_94_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_94, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_94);
	input_row_95_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_95, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_95);
	input_row_96_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_96, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_96);
	input_row_97_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_97, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_97);
	input_row_98_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_98, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_98);
	input_row_99_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_99, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_99);
	input_row_100_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_100, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_100);
	input_row_101_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_101, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_101);
	input_row_102_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_102, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_102);
	input_row_103_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_103, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_103);
	input_row_104_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_104, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_104);
	input_row_105_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_105, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_105);
	input_row_106_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_106, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_106);
	input_row_107_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_107, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_107);
	input_row_108_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_108, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_108);
	input_row_109_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_109, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_109);
	input_row_110_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_110, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_110);
	input_row_111_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_111, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_111);
	input_row_112_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_112, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_112);
	input_row_113_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_113, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_113);
	input_row_114_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_114, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_114);
	input_row_115_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_115, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_115);
	input_row_116_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_116, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_116);
	input_row_117_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_117, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_117);
	input_row_118_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_118, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_118);
	input_row_119_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_119, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_119);
	input_row_120_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_120, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_120);
	input_row_121_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_121, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_121);
	input_row_122_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_122, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_122);
	input_row_123_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_123, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_123);
	input_row_124_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_124, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_124);
	input_row_125_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_125, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_125);
	input_row_126_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_126, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_126);
	input_row_127_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_127, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_127);
	input_col_0_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_0, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_0);

	input_col_1_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_1, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_1);

	input_col_2_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_2, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_2);

	input_col_3_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_3, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_3);

	input_col_4_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_4, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_4);

	input_col_5_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_5, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_5);

	input_col_6_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_6, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_6);

	input_col_7_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_7, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_7);

	input_col_8_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_8, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_8);

	input_col_9_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_9, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_9);

	input_col_10_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_10, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_10);

	input_col_11_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_11, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_11);

	input_col_12_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_12, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_12);

	input_col_13_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_13, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_13);

	input_col_14_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_14, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_14);

	input_col_15_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_15, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_15);

	input_col_16_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_16, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_16);

	input_col_17_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_17, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_17);

	input_col_18_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_18, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_18);

	input_col_19_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_19, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_19);

	input_col_20_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_20, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_20);

	input_col_21_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_21, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_21);

	input_col_22_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_22, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_22);

	input_col_23_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_23, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_23);

	input_col_24_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_24, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_24);

	input_col_25_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_25, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_25);

	input_col_26_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_26, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_26);

	input_col_27_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_27, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_27);

	input_col_28_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_28, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_28);

	input_col_29_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_29, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_29);

	input_col_30_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_30, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_30);

	input_col_31_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_31, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_31);

	enable_ff_in: ff PORT MAP(D=>ENABLE, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>reg_ENABLE_in);
	sel_mux_reg: regnbit GENERIC MAP(N=>5) PORT MAP(D=>SEL_MUX, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>reg_SEL_MUX);

	MAC_0_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_0, data_out=>output_MAC_0_0);

	MAC_0_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_1, data_out=>output_MAC_0_1);

	MAC_0_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_2, data_out=>output_MAC_0_2);

	MAC_0_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_3, data_out=>output_MAC_0_3);

	MAC_0_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_4, data_out=>output_MAC_0_4);

	MAC_0_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_5, data_out=>output_MAC_0_5);

	MAC_0_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_6, data_out=>output_MAC_0_6);

	MAC_0_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_7, data_out=>output_MAC_0_7);

	MAC_0_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_8, data_out=>output_MAC_0_8);

	MAC_0_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_9, data_out=>output_MAC_0_9);

	MAC_0_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_10, data_out=>output_MAC_0_10);

	MAC_0_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_11, data_out=>output_MAC_0_11);

	MAC_0_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_12, data_out=>output_MAC_0_12);

	MAC_0_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_13, data_out=>output_MAC_0_13);

	MAC_0_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_14, data_out=>output_MAC_0_14);

	MAC_0_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_15, data_out=>output_MAC_0_15);

	MAC_0_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_16, data_out=>output_MAC_0_16);

	MAC_0_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_17, data_out=>output_MAC_0_17);

	MAC_0_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_18, data_out=>output_MAC_0_18);

	MAC_0_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_19, data_out=>output_MAC_0_19);

	MAC_0_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_20, data_out=>output_MAC_0_20);

	MAC_0_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_21, data_out=>output_MAC_0_21);

	MAC_0_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_22, data_out=>output_MAC_0_22);

	MAC_0_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_23, data_out=>output_MAC_0_23);

	MAC_0_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_24, data_out=>output_MAC_0_24);

	MAC_0_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_25, data_out=>output_MAC_0_25);

	MAC_0_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_26, data_out=>output_MAC_0_26);

	MAC_0_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_27, data_out=>output_MAC_0_27);

	MAC_0_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_28, data_out=>output_MAC_0_28);

	MAC_0_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_29, data_out=>output_MAC_0_29);

	MAC_0_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_30, data_out=>output_MAC_0_30);

	MAC_0_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_31, data_out=>output_MAC_0_31);

	MAC_1_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_0, data_out=>output_MAC_1_0);

	MAC_1_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_1, data_out=>output_MAC_1_1);

	MAC_1_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_2, data_out=>output_MAC_1_2);

	MAC_1_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_3, data_out=>output_MAC_1_3);

	MAC_1_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_4, data_out=>output_MAC_1_4);

	MAC_1_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_5, data_out=>output_MAC_1_5);

	MAC_1_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_6, data_out=>output_MAC_1_6);

	MAC_1_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_7, data_out=>output_MAC_1_7);

	MAC_1_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_8, data_out=>output_MAC_1_8);

	MAC_1_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_9, data_out=>output_MAC_1_9);

	MAC_1_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_10, data_out=>output_MAC_1_10);

	MAC_1_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_11, data_out=>output_MAC_1_11);

	MAC_1_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_12, data_out=>output_MAC_1_12);

	MAC_1_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_13, data_out=>output_MAC_1_13);

	MAC_1_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_14, data_out=>output_MAC_1_14);

	MAC_1_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_15, data_out=>output_MAC_1_15);

	MAC_1_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_16, data_out=>output_MAC_1_16);

	MAC_1_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_17, data_out=>output_MAC_1_17);

	MAC_1_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_18, data_out=>output_MAC_1_18);

	MAC_1_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_19, data_out=>output_MAC_1_19);

	MAC_1_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_20, data_out=>output_MAC_1_20);

	MAC_1_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_21, data_out=>output_MAC_1_21);

	MAC_1_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_22, data_out=>output_MAC_1_22);

	MAC_1_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_23, data_out=>output_MAC_1_23);

	MAC_1_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_24, data_out=>output_MAC_1_24);

	MAC_1_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_25, data_out=>output_MAC_1_25);

	MAC_1_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_26, data_out=>output_MAC_1_26);

	MAC_1_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_27, data_out=>output_MAC_1_27);

	MAC_1_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_28, data_out=>output_MAC_1_28);

	MAC_1_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_29, data_out=>output_MAC_1_29);

	MAC_1_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_30, data_out=>output_MAC_1_30);

	MAC_1_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_31, data_out=>output_MAC_1_31);

	MAC_2_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_0, data_out=>output_MAC_2_0);

	MAC_2_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_1, data_out=>output_MAC_2_1);

	MAC_2_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_2, data_out=>output_MAC_2_2);

	MAC_2_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_3, data_out=>output_MAC_2_3);

	MAC_2_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_4, data_out=>output_MAC_2_4);

	MAC_2_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_5, data_out=>output_MAC_2_5);

	MAC_2_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_6, data_out=>output_MAC_2_6);

	MAC_2_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_7, data_out=>output_MAC_2_7);

	MAC_2_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_8, data_out=>output_MAC_2_8);

	MAC_2_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_9, data_out=>output_MAC_2_9);

	MAC_2_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_10, data_out=>output_MAC_2_10);

	MAC_2_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_11, data_out=>output_MAC_2_11);

	MAC_2_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_12, data_out=>output_MAC_2_12);

	MAC_2_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_13, data_out=>output_MAC_2_13);

	MAC_2_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_14, data_out=>output_MAC_2_14);

	MAC_2_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_15, data_out=>output_MAC_2_15);

	MAC_2_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_16, data_out=>output_MAC_2_16);

	MAC_2_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_17, data_out=>output_MAC_2_17);

	MAC_2_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_18, data_out=>output_MAC_2_18);

	MAC_2_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_19, data_out=>output_MAC_2_19);

	MAC_2_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_20, data_out=>output_MAC_2_20);

	MAC_2_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_21, data_out=>output_MAC_2_21);

	MAC_2_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_22, data_out=>output_MAC_2_22);

	MAC_2_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_23, data_out=>output_MAC_2_23);

	MAC_2_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_24, data_out=>output_MAC_2_24);

	MAC_2_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_25, data_out=>output_MAC_2_25);

	MAC_2_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_26, data_out=>output_MAC_2_26);

	MAC_2_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_27, data_out=>output_MAC_2_27);

	MAC_2_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_28, data_out=>output_MAC_2_28);

	MAC_2_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_29, data_out=>output_MAC_2_29);

	MAC_2_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_30, data_out=>output_MAC_2_30);

	MAC_2_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_31, data_out=>output_MAC_2_31);

	MAC_3_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_0, data_out=>output_MAC_3_0);

	MAC_3_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_1, data_out=>output_MAC_3_1);

	MAC_3_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_2, data_out=>output_MAC_3_2);

	MAC_3_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_3, data_out=>output_MAC_3_3);

	MAC_3_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_4, data_out=>output_MAC_3_4);

	MAC_3_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_5, data_out=>output_MAC_3_5);

	MAC_3_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_6, data_out=>output_MAC_3_6);

	MAC_3_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_7, data_out=>output_MAC_3_7);

	MAC_3_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_8, data_out=>output_MAC_3_8);

	MAC_3_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_9, data_out=>output_MAC_3_9);

	MAC_3_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_10, data_out=>output_MAC_3_10);

	MAC_3_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_11, data_out=>output_MAC_3_11);

	MAC_3_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_12, data_out=>output_MAC_3_12);

	MAC_3_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_13, data_out=>output_MAC_3_13);

	MAC_3_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_14, data_out=>output_MAC_3_14);

	MAC_3_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_15, data_out=>output_MAC_3_15);

	MAC_3_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_16, data_out=>output_MAC_3_16);

	MAC_3_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_17, data_out=>output_MAC_3_17);

	MAC_3_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_18, data_out=>output_MAC_3_18);

	MAC_3_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_19, data_out=>output_MAC_3_19);

	MAC_3_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_20, data_out=>output_MAC_3_20);

	MAC_3_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_21, data_out=>output_MAC_3_21);

	MAC_3_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_22, data_out=>output_MAC_3_22);

	MAC_3_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_23, data_out=>output_MAC_3_23);

	MAC_3_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_24, data_out=>output_MAC_3_24);

	MAC_3_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_25, data_out=>output_MAC_3_25);

	MAC_3_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_26, data_out=>output_MAC_3_26);

	MAC_3_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_27, data_out=>output_MAC_3_27);

	MAC_3_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_28, data_out=>output_MAC_3_28);

	MAC_3_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_29, data_out=>output_MAC_3_29);

	MAC_3_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_30, data_out=>output_MAC_3_30);

	MAC_3_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_31, data_out=>output_MAC_3_31);

	MAC_4_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_0, data_out=>output_MAC_4_0);

	MAC_4_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_1, data_out=>output_MAC_4_1);

	MAC_4_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_2, data_out=>output_MAC_4_2);

	MAC_4_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_3, data_out=>output_MAC_4_3);

	MAC_4_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_4, data_out=>output_MAC_4_4);

	MAC_4_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_5, data_out=>output_MAC_4_5);

	MAC_4_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_6, data_out=>output_MAC_4_6);

	MAC_4_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_7, data_out=>output_MAC_4_7);

	MAC_4_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_8, data_out=>output_MAC_4_8);

	MAC_4_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_9, data_out=>output_MAC_4_9);

	MAC_4_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_10, data_out=>output_MAC_4_10);

	MAC_4_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_11, data_out=>output_MAC_4_11);

	MAC_4_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_12, data_out=>output_MAC_4_12);

	MAC_4_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_13, data_out=>output_MAC_4_13);

	MAC_4_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_14, data_out=>output_MAC_4_14);

	MAC_4_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_15, data_out=>output_MAC_4_15);

	MAC_4_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_16, data_out=>output_MAC_4_16);

	MAC_4_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_17, data_out=>output_MAC_4_17);

	MAC_4_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_18, data_out=>output_MAC_4_18);

	MAC_4_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_19, data_out=>output_MAC_4_19);

	MAC_4_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_20, data_out=>output_MAC_4_20);

	MAC_4_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_21, data_out=>output_MAC_4_21);

	MAC_4_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_22, data_out=>output_MAC_4_22);

	MAC_4_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_23, data_out=>output_MAC_4_23);

	MAC_4_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_24, data_out=>output_MAC_4_24);

	MAC_4_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_25, data_out=>output_MAC_4_25);

	MAC_4_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_26, data_out=>output_MAC_4_26);

	MAC_4_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_27, data_out=>output_MAC_4_27);

	MAC_4_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_28, data_out=>output_MAC_4_28);

	MAC_4_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_29, data_out=>output_MAC_4_29);

	MAC_4_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_30, data_out=>output_MAC_4_30);

	MAC_4_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_31, data_out=>output_MAC_4_31);

	MAC_5_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_0, data_out=>output_MAC_5_0);

	MAC_5_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_1, data_out=>output_MAC_5_1);

	MAC_5_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_2, data_out=>output_MAC_5_2);

	MAC_5_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_3, data_out=>output_MAC_5_3);

	MAC_5_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_4, data_out=>output_MAC_5_4);

	MAC_5_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_5, data_out=>output_MAC_5_5);

	MAC_5_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_6, data_out=>output_MAC_5_6);

	MAC_5_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_7, data_out=>output_MAC_5_7);

	MAC_5_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_8, data_out=>output_MAC_5_8);

	MAC_5_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_9, data_out=>output_MAC_5_9);

	MAC_5_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_10, data_out=>output_MAC_5_10);

	MAC_5_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_11, data_out=>output_MAC_5_11);

	MAC_5_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_12, data_out=>output_MAC_5_12);

	MAC_5_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_13, data_out=>output_MAC_5_13);

	MAC_5_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_14, data_out=>output_MAC_5_14);

	MAC_5_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_15, data_out=>output_MAC_5_15);

	MAC_5_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_16, data_out=>output_MAC_5_16);

	MAC_5_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_17, data_out=>output_MAC_5_17);

	MAC_5_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_18, data_out=>output_MAC_5_18);

	MAC_5_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_19, data_out=>output_MAC_5_19);

	MAC_5_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_20, data_out=>output_MAC_5_20);

	MAC_5_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_21, data_out=>output_MAC_5_21);

	MAC_5_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_22, data_out=>output_MAC_5_22);

	MAC_5_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_23, data_out=>output_MAC_5_23);

	MAC_5_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_24, data_out=>output_MAC_5_24);

	MAC_5_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_25, data_out=>output_MAC_5_25);

	MAC_5_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_26, data_out=>output_MAC_5_26);

	MAC_5_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_27, data_out=>output_MAC_5_27);

	MAC_5_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_28, data_out=>output_MAC_5_28);

	MAC_5_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_29, data_out=>output_MAC_5_29);

	MAC_5_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_30, data_out=>output_MAC_5_30);

	MAC_5_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_31, data_out=>output_MAC_5_31);

	MAC_6_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_0, data_out=>output_MAC_6_0);

	MAC_6_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_1, data_out=>output_MAC_6_1);

	MAC_6_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_2, data_out=>output_MAC_6_2);

	MAC_6_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_3, data_out=>output_MAC_6_3);

	MAC_6_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_4, data_out=>output_MAC_6_4);

	MAC_6_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_5, data_out=>output_MAC_6_5);

	MAC_6_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_6, data_out=>output_MAC_6_6);

	MAC_6_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_7, data_out=>output_MAC_6_7);

	MAC_6_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_8, data_out=>output_MAC_6_8);

	MAC_6_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_9, data_out=>output_MAC_6_9);

	MAC_6_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_10, data_out=>output_MAC_6_10);

	MAC_6_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_11, data_out=>output_MAC_6_11);

	MAC_6_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_12, data_out=>output_MAC_6_12);

	MAC_6_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_13, data_out=>output_MAC_6_13);

	MAC_6_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_14, data_out=>output_MAC_6_14);

	MAC_6_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_15, data_out=>output_MAC_6_15);

	MAC_6_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_16, data_out=>output_MAC_6_16);

	MAC_6_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_17, data_out=>output_MAC_6_17);

	MAC_6_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_18, data_out=>output_MAC_6_18);

	MAC_6_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_19, data_out=>output_MAC_6_19);

	MAC_6_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_20, data_out=>output_MAC_6_20);

	MAC_6_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_21, data_out=>output_MAC_6_21);

	MAC_6_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_22, data_out=>output_MAC_6_22);

	MAC_6_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_23, data_out=>output_MAC_6_23);

	MAC_6_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_24, data_out=>output_MAC_6_24);

	MAC_6_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_25, data_out=>output_MAC_6_25);

	MAC_6_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_26, data_out=>output_MAC_6_26);

	MAC_6_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_27, data_out=>output_MAC_6_27);

	MAC_6_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_28, data_out=>output_MAC_6_28);

	MAC_6_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_29, data_out=>output_MAC_6_29);

	MAC_6_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_30, data_out=>output_MAC_6_30);

	MAC_6_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_31, data_out=>output_MAC_6_31);

	MAC_7_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_0, data_out=>output_MAC_7_0);

	MAC_7_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_1, data_out=>output_MAC_7_1);

	MAC_7_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_2, data_out=>output_MAC_7_2);

	MAC_7_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_3, data_out=>output_MAC_7_3);

	MAC_7_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_4, data_out=>output_MAC_7_4);

	MAC_7_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_5, data_out=>output_MAC_7_5);

	MAC_7_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_6, data_out=>output_MAC_7_6);

	MAC_7_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_7, data_out=>output_MAC_7_7);

	MAC_7_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_8, data_out=>output_MAC_7_8);

	MAC_7_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_9, data_out=>output_MAC_7_9);

	MAC_7_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_10, data_out=>output_MAC_7_10);

	MAC_7_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_11, data_out=>output_MAC_7_11);

	MAC_7_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_12, data_out=>output_MAC_7_12);

	MAC_7_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_13, data_out=>output_MAC_7_13);

	MAC_7_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_14, data_out=>output_MAC_7_14);

	MAC_7_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_15, data_out=>output_MAC_7_15);

	MAC_7_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_16, data_out=>output_MAC_7_16);

	MAC_7_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_17, data_out=>output_MAC_7_17);

	MAC_7_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_18, data_out=>output_MAC_7_18);

	MAC_7_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_19, data_out=>output_MAC_7_19);

	MAC_7_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_20, data_out=>output_MAC_7_20);

	MAC_7_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_21, data_out=>output_MAC_7_21);

	MAC_7_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_22, data_out=>output_MAC_7_22);

	MAC_7_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_23, data_out=>output_MAC_7_23);

	MAC_7_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_24, data_out=>output_MAC_7_24);

	MAC_7_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_25, data_out=>output_MAC_7_25);

	MAC_7_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_26, data_out=>output_MAC_7_26);

	MAC_7_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_27, data_out=>output_MAC_7_27);

	MAC_7_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_28, data_out=>output_MAC_7_28);

	MAC_7_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_29, data_out=>output_MAC_7_29);

	MAC_7_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_30, data_out=>output_MAC_7_30);

	MAC_7_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_31, data_out=>output_MAC_7_31);

	MAC_8_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_0, data_out=>output_MAC_8_0);

	MAC_8_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_1, data_out=>output_MAC_8_1);

	MAC_8_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_2, data_out=>output_MAC_8_2);

	MAC_8_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_3, data_out=>output_MAC_8_3);

	MAC_8_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_4, data_out=>output_MAC_8_4);

	MAC_8_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_5, data_out=>output_MAC_8_5);

	MAC_8_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_6, data_out=>output_MAC_8_6);

	MAC_8_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_7, data_out=>output_MAC_8_7);

	MAC_8_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_8, data_out=>output_MAC_8_8);

	MAC_8_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_9, data_out=>output_MAC_8_9);

	MAC_8_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_10, data_out=>output_MAC_8_10);

	MAC_8_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_11, data_out=>output_MAC_8_11);

	MAC_8_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_12, data_out=>output_MAC_8_12);

	MAC_8_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_13, data_out=>output_MAC_8_13);

	MAC_8_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_14, data_out=>output_MAC_8_14);

	MAC_8_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_15, data_out=>output_MAC_8_15);

	MAC_8_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_16, data_out=>output_MAC_8_16);

	MAC_8_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_17, data_out=>output_MAC_8_17);

	MAC_8_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_18, data_out=>output_MAC_8_18);

	MAC_8_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_19, data_out=>output_MAC_8_19);

	MAC_8_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_20, data_out=>output_MAC_8_20);

	MAC_8_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_21, data_out=>output_MAC_8_21);

	MAC_8_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_22, data_out=>output_MAC_8_22);

	MAC_8_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_23, data_out=>output_MAC_8_23);

	MAC_8_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_24, data_out=>output_MAC_8_24);

	MAC_8_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_25, data_out=>output_MAC_8_25);

	MAC_8_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_26, data_out=>output_MAC_8_26);

	MAC_8_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_27, data_out=>output_MAC_8_27);

	MAC_8_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_28, data_out=>output_MAC_8_28);

	MAC_8_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_29, data_out=>output_MAC_8_29);

	MAC_8_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_30, data_out=>output_MAC_8_30);

	MAC_8_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_31, data_out=>output_MAC_8_31);

	MAC_9_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_0, data_out=>output_MAC_9_0);

	MAC_9_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_1, data_out=>output_MAC_9_1);

	MAC_9_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_2, data_out=>output_MAC_9_2);

	MAC_9_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_3, data_out=>output_MAC_9_3);

	MAC_9_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_4, data_out=>output_MAC_9_4);

	MAC_9_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_5, data_out=>output_MAC_9_5);

	MAC_9_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_6, data_out=>output_MAC_9_6);

	MAC_9_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_7, data_out=>output_MAC_9_7);

	MAC_9_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_8, data_out=>output_MAC_9_8);

	MAC_9_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_9, data_out=>output_MAC_9_9);

	MAC_9_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_10, data_out=>output_MAC_9_10);

	MAC_9_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_11, data_out=>output_MAC_9_11);

	MAC_9_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_12, data_out=>output_MAC_9_12);

	MAC_9_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_13, data_out=>output_MAC_9_13);

	MAC_9_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_14, data_out=>output_MAC_9_14);

	MAC_9_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_15, data_out=>output_MAC_9_15);

	MAC_9_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_16, data_out=>output_MAC_9_16);

	MAC_9_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_17, data_out=>output_MAC_9_17);

	MAC_9_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_18, data_out=>output_MAC_9_18);

	MAC_9_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_19, data_out=>output_MAC_9_19);

	MAC_9_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_20, data_out=>output_MAC_9_20);

	MAC_9_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_21, data_out=>output_MAC_9_21);

	MAC_9_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_22, data_out=>output_MAC_9_22);

	MAC_9_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_23, data_out=>output_MAC_9_23);

	MAC_9_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_24, data_out=>output_MAC_9_24);

	MAC_9_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_25, data_out=>output_MAC_9_25);

	MAC_9_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_26, data_out=>output_MAC_9_26);

	MAC_9_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_27, data_out=>output_MAC_9_27);

	MAC_9_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_28, data_out=>output_MAC_9_28);

	MAC_9_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_29, data_out=>output_MAC_9_29);

	MAC_9_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_30, data_out=>output_MAC_9_30);

	MAC_9_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_31, data_out=>output_MAC_9_31);

	MAC_10_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_0, data_out=>output_MAC_10_0);

	MAC_10_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_1, data_out=>output_MAC_10_1);

	MAC_10_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_2, data_out=>output_MAC_10_2);

	MAC_10_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_3, data_out=>output_MAC_10_3);

	MAC_10_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_4, data_out=>output_MAC_10_4);

	MAC_10_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_5, data_out=>output_MAC_10_5);

	MAC_10_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_6, data_out=>output_MAC_10_6);

	MAC_10_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_7, data_out=>output_MAC_10_7);

	MAC_10_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_8, data_out=>output_MAC_10_8);

	MAC_10_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_9, data_out=>output_MAC_10_9);

	MAC_10_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_10, data_out=>output_MAC_10_10);

	MAC_10_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_11, data_out=>output_MAC_10_11);

	MAC_10_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_12, data_out=>output_MAC_10_12);

	MAC_10_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_13, data_out=>output_MAC_10_13);

	MAC_10_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_14, data_out=>output_MAC_10_14);

	MAC_10_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_15, data_out=>output_MAC_10_15);

	MAC_10_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_16, data_out=>output_MAC_10_16);

	MAC_10_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_17, data_out=>output_MAC_10_17);

	MAC_10_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_18, data_out=>output_MAC_10_18);

	MAC_10_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_19, data_out=>output_MAC_10_19);

	MAC_10_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_20, data_out=>output_MAC_10_20);

	MAC_10_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_21, data_out=>output_MAC_10_21);

	MAC_10_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_22, data_out=>output_MAC_10_22);

	MAC_10_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_23, data_out=>output_MAC_10_23);

	MAC_10_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_24, data_out=>output_MAC_10_24);

	MAC_10_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_25, data_out=>output_MAC_10_25);

	MAC_10_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_26, data_out=>output_MAC_10_26);

	MAC_10_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_27, data_out=>output_MAC_10_27);

	MAC_10_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_28, data_out=>output_MAC_10_28);

	MAC_10_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_29, data_out=>output_MAC_10_29);

	MAC_10_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_30, data_out=>output_MAC_10_30);

	MAC_10_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_31, data_out=>output_MAC_10_31);

	MAC_11_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_0, data_out=>output_MAC_11_0);

	MAC_11_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_1, data_out=>output_MAC_11_1);

	MAC_11_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_2, data_out=>output_MAC_11_2);

	MAC_11_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_3, data_out=>output_MAC_11_3);

	MAC_11_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_4, data_out=>output_MAC_11_4);

	MAC_11_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_5, data_out=>output_MAC_11_5);

	MAC_11_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_6, data_out=>output_MAC_11_6);

	MAC_11_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_7, data_out=>output_MAC_11_7);

	MAC_11_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_8, data_out=>output_MAC_11_8);

	MAC_11_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_9, data_out=>output_MAC_11_9);

	MAC_11_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_10, data_out=>output_MAC_11_10);

	MAC_11_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_11, data_out=>output_MAC_11_11);

	MAC_11_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_12, data_out=>output_MAC_11_12);

	MAC_11_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_13, data_out=>output_MAC_11_13);

	MAC_11_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_14, data_out=>output_MAC_11_14);

	MAC_11_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_15, data_out=>output_MAC_11_15);

	MAC_11_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_16, data_out=>output_MAC_11_16);

	MAC_11_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_17, data_out=>output_MAC_11_17);

	MAC_11_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_18, data_out=>output_MAC_11_18);

	MAC_11_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_19, data_out=>output_MAC_11_19);

	MAC_11_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_20, data_out=>output_MAC_11_20);

	MAC_11_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_21, data_out=>output_MAC_11_21);

	MAC_11_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_22, data_out=>output_MAC_11_22);

	MAC_11_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_23, data_out=>output_MAC_11_23);

	MAC_11_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_24, data_out=>output_MAC_11_24);

	MAC_11_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_25, data_out=>output_MAC_11_25);

	MAC_11_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_26, data_out=>output_MAC_11_26);

	MAC_11_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_27, data_out=>output_MAC_11_27);

	MAC_11_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_28, data_out=>output_MAC_11_28);

	MAC_11_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_29, data_out=>output_MAC_11_29);

	MAC_11_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_30, data_out=>output_MAC_11_30);

	MAC_11_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_31, data_out=>output_MAC_11_31);

	MAC_12_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_0, data_out=>output_MAC_12_0);

	MAC_12_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_1, data_out=>output_MAC_12_1);

	MAC_12_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_2, data_out=>output_MAC_12_2);

	MAC_12_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_3, data_out=>output_MAC_12_3);

	MAC_12_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_4, data_out=>output_MAC_12_4);

	MAC_12_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_5, data_out=>output_MAC_12_5);

	MAC_12_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_6, data_out=>output_MAC_12_6);

	MAC_12_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_7, data_out=>output_MAC_12_7);

	MAC_12_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_8, data_out=>output_MAC_12_8);

	MAC_12_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_9, data_out=>output_MAC_12_9);

	MAC_12_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_10, data_out=>output_MAC_12_10);

	MAC_12_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_11, data_out=>output_MAC_12_11);

	MAC_12_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_12, data_out=>output_MAC_12_12);

	MAC_12_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_13, data_out=>output_MAC_12_13);

	MAC_12_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_14, data_out=>output_MAC_12_14);

	MAC_12_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_15, data_out=>output_MAC_12_15);

	MAC_12_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_16, data_out=>output_MAC_12_16);

	MAC_12_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_17, data_out=>output_MAC_12_17);

	MAC_12_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_18, data_out=>output_MAC_12_18);

	MAC_12_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_19, data_out=>output_MAC_12_19);

	MAC_12_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_20, data_out=>output_MAC_12_20);

	MAC_12_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_21, data_out=>output_MAC_12_21);

	MAC_12_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_22, data_out=>output_MAC_12_22);

	MAC_12_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_23, data_out=>output_MAC_12_23);

	MAC_12_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_24, data_out=>output_MAC_12_24);

	MAC_12_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_25, data_out=>output_MAC_12_25);

	MAC_12_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_26, data_out=>output_MAC_12_26);

	MAC_12_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_27, data_out=>output_MAC_12_27);

	MAC_12_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_28, data_out=>output_MAC_12_28);

	MAC_12_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_29, data_out=>output_MAC_12_29);

	MAC_12_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_30, data_out=>output_MAC_12_30);

	MAC_12_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_31, data_out=>output_MAC_12_31);

	MAC_13_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_0, data_out=>output_MAC_13_0);

	MAC_13_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_1, data_out=>output_MAC_13_1);

	MAC_13_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_2, data_out=>output_MAC_13_2);

	MAC_13_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_3, data_out=>output_MAC_13_3);

	MAC_13_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_4, data_out=>output_MAC_13_4);

	MAC_13_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_5, data_out=>output_MAC_13_5);

	MAC_13_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_6, data_out=>output_MAC_13_6);

	MAC_13_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_7, data_out=>output_MAC_13_7);

	MAC_13_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_8, data_out=>output_MAC_13_8);

	MAC_13_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_9, data_out=>output_MAC_13_9);

	MAC_13_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_10, data_out=>output_MAC_13_10);

	MAC_13_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_11, data_out=>output_MAC_13_11);

	MAC_13_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_12, data_out=>output_MAC_13_12);

	MAC_13_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_13, data_out=>output_MAC_13_13);

	MAC_13_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_14, data_out=>output_MAC_13_14);

	MAC_13_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_15, data_out=>output_MAC_13_15);

	MAC_13_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_16, data_out=>output_MAC_13_16);

	MAC_13_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_17, data_out=>output_MAC_13_17);

	MAC_13_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_18, data_out=>output_MAC_13_18);

	MAC_13_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_19, data_out=>output_MAC_13_19);

	MAC_13_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_20, data_out=>output_MAC_13_20);

	MAC_13_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_21, data_out=>output_MAC_13_21);

	MAC_13_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_22, data_out=>output_MAC_13_22);

	MAC_13_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_23, data_out=>output_MAC_13_23);

	MAC_13_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_24, data_out=>output_MAC_13_24);

	MAC_13_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_25, data_out=>output_MAC_13_25);

	MAC_13_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_26, data_out=>output_MAC_13_26);

	MAC_13_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_27, data_out=>output_MAC_13_27);

	MAC_13_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_28, data_out=>output_MAC_13_28);

	MAC_13_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_29, data_out=>output_MAC_13_29);

	MAC_13_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_30, data_out=>output_MAC_13_30);

	MAC_13_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_31, data_out=>output_MAC_13_31);

	MAC_14_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_0, data_out=>output_MAC_14_0);

	MAC_14_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_1, data_out=>output_MAC_14_1);

	MAC_14_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_2, data_out=>output_MAC_14_2);

	MAC_14_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_3, data_out=>output_MAC_14_3);

	MAC_14_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_4, data_out=>output_MAC_14_4);

	MAC_14_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_5, data_out=>output_MAC_14_5);

	MAC_14_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_6, data_out=>output_MAC_14_6);

	MAC_14_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_7, data_out=>output_MAC_14_7);

	MAC_14_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_8, data_out=>output_MAC_14_8);

	MAC_14_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_9, data_out=>output_MAC_14_9);

	MAC_14_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_10, data_out=>output_MAC_14_10);

	MAC_14_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_11, data_out=>output_MAC_14_11);

	MAC_14_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_12, data_out=>output_MAC_14_12);

	MAC_14_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_13, data_out=>output_MAC_14_13);

	MAC_14_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_14, data_out=>output_MAC_14_14);

	MAC_14_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_15, data_out=>output_MAC_14_15);

	MAC_14_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_16, data_out=>output_MAC_14_16);

	MAC_14_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_17, data_out=>output_MAC_14_17);

	MAC_14_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_18, data_out=>output_MAC_14_18);

	MAC_14_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_19, data_out=>output_MAC_14_19);

	MAC_14_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_20, data_out=>output_MAC_14_20);

	MAC_14_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_21, data_out=>output_MAC_14_21);

	MAC_14_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_22, data_out=>output_MAC_14_22);

	MAC_14_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_23, data_out=>output_MAC_14_23);

	MAC_14_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_24, data_out=>output_MAC_14_24);

	MAC_14_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_25, data_out=>output_MAC_14_25);

	MAC_14_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_26, data_out=>output_MAC_14_26);

	MAC_14_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_27, data_out=>output_MAC_14_27);

	MAC_14_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_28, data_out=>output_MAC_14_28);

	MAC_14_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_29, data_out=>output_MAC_14_29);

	MAC_14_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_30, data_out=>output_MAC_14_30);

	MAC_14_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_31, data_out=>output_MAC_14_31);

	MAC_15_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_0, data_out=>output_MAC_15_0);

	MAC_15_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_1, data_out=>output_MAC_15_1);

	MAC_15_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_2, data_out=>output_MAC_15_2);

	MAC_15_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_3, data_out=>output_MAC_15_3);

	MAC_15_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_4, data_out=>output_MAC_15_4);

	MAC_15_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_5, data_out=>output_MAC_15_5);

	MAC_15_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_6, data_out=>output_MAC_15_6);

	MAC_15_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_7, data_out=>output_MAC_15_7);

	MAC_15_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_8, data_out=>output_MAC_15_8);

	MAC_15_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_9, data_out=>output_MAC_15_9);

	MAC_15_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_10, data_out=>output_MAC_15_10);

	MAC_15_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_11, data_out=>output_MAC_15_11);

	MAC_15_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_12, data_out=>output_MAC_15_12);

	MAC_15_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_13, data_out=>output_MAC_15_13);

	MAC_15_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_14, data_out=>output_MAC_15_14);

	MAC_15_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_15, data_out=>output_MAC_15_15);

	MAC_15_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_16, data_out=>output_MAC_15_16);

	MAC_15_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_17, data_out=>output_MAC_15_17);

	MAC_15_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_18, data_out=>output_MAC_15_18);

	MAC_15_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_19, data_out=>output_MAC_15_19);

	MAC_15_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_20, data_out=>output_MAC_15_20);

	MAC_15_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_21, data_out=>output_MAC_15_21);

	MAC_15_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_22, data_out=>output_MAC_15_22);

	MAC_15_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_23, data_out=>output_MAC_15_23);

	MAC_15_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_24, data_out=>output_MAC_15_24);

	MAC_15_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_25, data_out=>output_MAC_15_25);

	MAC_15_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_26, data_out=>output_MAC_15_26);

	MAC_15_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_27, data_out=>output_MAC_15_27);

	MAC_15_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_28, data_out=>output_MAC_15_28);

	MAC_15_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_29, data_out=>output_MAC_15_29);

	MAC_15_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_30, data_out=>output_MAC_15_30);

	MAC_15_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_31, data_out=>output_MAC_15_31);

	MAC_16_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_0, data_out=>output_MAC_16_0);

	MAC_16_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_1, data_out=>output_MAC_16_1);

	MAC_16_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_2, data_out=>output_MAC_16_2);

	MAC_16_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_3, data_out=>output_MAC_16_3);

	MAC_16_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_4, data_out=>output_MAC_16_4);

	MAC_16_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_5, data_out=>output_MAC_16_5);

	MAC_16_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_6, data_out=>output_MAC_16_6);

	MAC_16_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_7, data_out=>output_MAC_16_7);

	MAC_16_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_8, data_out=>output_MAC_16_8);

	MAC_16_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_9, data_out=>output_MAC_16_9);

	MAC_16_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_10, data_out=>output_MAC_16_10);

	MAC_16_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_11, data_out=>output_MAC_16_11);

	MAC_16_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_12, data_out=>output_MAC_16_12);

	MAC_16_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_13, data_out=>output_MAC_16_13);

	MAC_16_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_14, data_out=>output_MAC_16_14);

	MAC_16_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_15, data_out=>output_MAC_16_15);

	MAC_16_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_16, data_out=>output_MAC_16_16);

	MAC_16_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_17, data_out=>output_MAC_16_17);

	MAC_16_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_18, data_out=>output_MAC_16_18);

	MAC_16_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_19, data_out=>output_MAC_16_19);

	MAC_16_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_20, data_out=>output_MAC_16_20);

	MAC_16_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_21, data_out=>output_MAC_16_21);

	MAC_16_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_22, data_out=>output_MAC_16_22);

	MAC_16_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_23, data_out=>output_MAC_16_23);

	MAC_16_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_24, data_out=>output_MAC_16_24);

	MAC_16_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_25, data_out=>output_MAC_16_25);

	MAC_16_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_26, data_out=>output_MAC_16_26);

	MAC_16_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_27, data_out=>output_MAC_16_27);

	MAC_16_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_28, data_out=>output_MAC_16_28);

	MAC_16_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_29, data_out=>output_MAC_16_29);

	MAC_16_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_30, data_out=>output_MAC_16_30);

	MAC_16_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_31, data_out=>output_MAC_16_31);

	MAC_17_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_0, data_out=>output_MAC_17_0);

	MAC_17_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_1, data_out=>output_MAC_17_1);

	MAC_17_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_2, data_out=>output_MAC_17_2);

	MAC_17_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_3, data_out=>output_MAC_17_3);

	MAC_17_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_4, data_out=>output_MAC_17_4);

	MAC_17_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_5, data_out=>output_MAC_17_5);

	MAC_17_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_6, data_out=>output_MAC_17_6);

	MAC_17_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_7, data_out=>output_MAC_17_7);

	MAC_17_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_8, data_out=>output_MAC_17_8);

	MAC_17_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_9, data_out=>output_MAC_17_9);

	MAC_17_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_10, data_out=>output_MAC_17_10);

	MAC_17_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_11, data_out=>output_MAC_17_11);

	MAC_17_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_12, data_out=>output_MAC_17_12);

	MAC_17_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_13, data_out=>output_MAC_17_13);

	MAC_17_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_14, data_out=>output_MAC_17_14);

	MAC_17_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_15, data_out=>output_MAC_17_15);

	MAC_17_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_16, data_out=>output_MAC_17_16);

	MAC_17_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_17, data_out=>output_MAC_17_17);

	MAC_17_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_18, data_out=>output_MAC_17_18);

	MAC_17_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_19, data_out=>output_MAC_17_19);

	MAC_17_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_20, data_out=>output_MAC_17_20);

	MAC_17_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_21, data_out=>output_MAC_17_21);

	MAC_17_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_22, data_out=>output_MAC_17_22);

	MAC_17_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_23, data_out=>output_MAC_17_23);

	MAC_17_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_24, data_out=>output_MAC_17_24);

	MAC_17_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_25, data_out=>output_MAC_17_25);

	MAC_17_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_26, data_out=>output_MAC_17_26);

	MAC_17_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_27, data_out=>output_MAC_17_27);

	MAC_17_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_28, data_out=>output_MAC_17_28);

	MAC_17_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_29, data_out=>output_MAC_17_29);

	MAC_17_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_30, data_out=>output_MAC_17_30);

	MAC_17_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_31, data_out=>output_MAC_17_31);

	MAC_18_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_0, data_out=>output_MAC_18_0);

	MAC_18_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_1, data_out=>output_MAC_18_1);

	MAC_18_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_2, data_out=>output_MAC_18_2);

	MAC_18_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_3, data_out=>output_MAC_18_3);

	MAC_18_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_4, data_out=>output_MAC_18_4);

	MAC_18_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_5, data_out=>output_MAC_18_5);

	MAC_18_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_6, data_out=>output_MAC_18_6);

	MAC_18_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_7, data_out=>output_MAC_18_7);

	MAC_18_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_8, data_out=>output_MAC_18_8);

	MAC_18_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_9, data_out=>output_MAC_18_9);

	MAC_18_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_10, data_out=>output_MAC_18_10);

	MAC_18_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_11, data_out=>output_MAC_18_11);

	MAC_18_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_12, data_out=>output_MAC_18_12);

	MAC_18_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_13, data_out=>output_MAC_18_13);

	MAC_18_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_14, data_out=>output_MAC_18_14);

	MAC_18_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_15, data_out=>output_MAC_18_15);

	MAC_18_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_16, data_out=>output_MAC_18_16);

	MAC_18_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_17, data_out=>output_MAC_18_17);

	MAC_18_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_18, data_out=>output_MAC_18_18);

	MAC_18_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_19, data_out=>output_MAC_18_19);

	MAC_18_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_20, data_out=>output_MAC_18_20);

	MAC_18_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_21, data_out=>output_MAC_18_21);

	MAC_18_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_22, data_out=>output_MAC_18_22);

	MAC_18_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_23, data_out=>output_MAC_18_23);

	MAC_18_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_24, data_out=>output_MAC_18_24);

	MAC_18_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_25, data_out=>output_MAC_18_25);

	MAC_18_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_26, data_out=>output_MAC_18_26);

	MAC_18_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_27, data_out=>output_MAC_18_27);

	MAC_18_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_28, data_out=>output_MAC_18_28);

	MAC_18_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_29, data_out=>output_MAC_18_29);

	MAC_18_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_30, data_out=>output_MAC_18_30);

	MAC_18_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_31, data_out=>output_MAC_18_31);

	MAC_19_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_0, data_out=>output_MAC_19_0);

	MAC_19_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_1, data_out=>output_MAC_19_1);

	MAC_19_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_2, data_out=>output_MAC_19_2);

	MAC_19_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_3, data_out=>output_MAC_19_3);

	MAC_19_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_4, data_out=>output_MAC_19_4);

	MAC_19_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_5, data_out=>output_MAC_19_5);

	MAC_19_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_6, data_out=>output_MAC_19_6);

	MAC_19_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_7, data_out=>output_MAC_19_7);

	MAC_19_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_8, data_out=>output_MAC_19_8);

	MAC_19_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_9, data_out=>output_MAC_19_9);

	MAC_19_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_10, data_out=>output_MAC_19_10);

	MAC_19_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_11, data_out=>output_MAC_19_11);

	MAC_19_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_12, data_out=>output_MAC_19_12);

	MAC_19_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_13, data_out=>output_MAC_19_13);

	MAC_19_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_14, data_out=>output_MAC_19_14);

	MAC_19_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_15, data_out=>output_MAC_19_15);

	MAC_19_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_16, data_out=>output_MAC_19_16);

	MAC_19_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_17, data_out=>output_MAC_19_17);

	MAC_19_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_18, data_out=>output_MAC_19_18);

	MAC_19_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_19, data_out=>output_MAC_19_19);

	MAC_19_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_20, data_out=>output_MAC_19_20);

	MAC_19_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_21, data_out=>output_MAC_19_21);

	MAC_19_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_22, data_out=>output_MAC_19_22);

	MAC_19_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_23, data_out=>output_MAC_19_23);

	MAC_19_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_24, data_out=>output_MAC_19_24);

	MAC_19_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_25, data_out=>output_MAC_19_25);

	MAC_19_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_26, data_out=>output_MAC_19_26);

	MAC_19_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_27, data_out=>output_MAC_19_27);

	MAC_19_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_28, data_out=>output_MAC_19_28);

	MAC_19_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_29, data_out=>output_MAC_19_29);

	MAC_19_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_30, data_out=>output_MAC_19_30);

	MAC_19_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_31, data_out=>output_MAC_19_31);

	MAC_20_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_0, data_out=>output_MAC_20_0);

	MAC_20_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_1, data_out=>output_MAC_20_1);

	MAC_20_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_2, data_out=>output_MAC_20_2);

	MAC_20_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_3, data_out=>output_MAC_20_3);

	MAC_20_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_4, data_out=>output_MAC_20_4);

	MAC_20_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_5, data_out=>output_MAC_20_5);

	MAC_20_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_6, data_out=>output_MAC_20_6);

	MAC_20_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_7, data_out=>output_MAC_20_7);

	MAC_20_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_8, data_out=>output_MAC_20_8);

	MAC_20_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_9, data_out=>output_MAC_20_9);

	MAC_20_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_10, data_out=>output_MAC_20_10);

	MAC_20_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_11, data_out=>output_MAC_20_11);

	MAC_20_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_12, data_out=>output_MAC_20_12);

	MAC_20_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_13, data_out=>output_MAC_20_13);

	MAC_20_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_14, data_out=>output_MAC_20_14);

	MAC_20_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_15, data_out=>output_MAC_20_15);

	MAC_20_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_16, data_out=>output_MAC_20_16);

	MAC_20_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_17, data_out=>output_MAC_20_17);

	MAC_20_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_18, data_out=>output_MAC_20_18);

	MAC_20_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_19, data_out=>output_MAC_20_19);

	MAC_20_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_20, data_out=>output_MAC_20_20);

	MAC_20_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_21, data_out=>output_MAC_20_21);

	MAC_20_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_22, data_out=>output_MAC_20_22);

	MAC_20_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_23, data_out=>output_MAC_20_23);

	MAC_20_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_24, data_out=>output_MAC_20_24);

	MAC_20_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_25, data_out=>output_MAC_20_25);

	MAC_20_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_26, data_out=>output_MAC_20_26);

	MAC_20_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_27, data_out=>output_MAC_20_27);

	MAC_20_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_28, data_out=>output_MAC_20_28);

	MAC_20_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_29, data_out=>output_MAC_20_29);

	MAC_20_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_30, data_out=>output_MAC_20_30);

	MAC_20_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_31, data_out=>output_MAC_20_31);

	MAC_21_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_0, data_out=>output_MAC_21_0);

	MAC_21_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_1, data_out=>output_MAC_21_1);

	MAC_21_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_2, data_out=>output_MAC_21_2);

	MAC_21_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_3, data_out=>output_MAC_21_3);

	MAC_21_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_4, data_out=>output_MAC_21_4);

	MAC_21_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_5, data_out=>output_MAC_21_5);

	MAC_21_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_6, data_out=>output_MAC_21_6);

	MAC_21_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_7, data_out=>output_MAC_21_7);

	MAC_21_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_8, data_out=>output_MAC_21_8);

	MAC_21_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_9, data_out=>output_MAC_21_9);

	MAC_21_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_10, data_out=>output_MAC_21_10);

	MAC_21_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_11, data_out=>output_MAC_21_11);

	MAC_21_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_12, data_out=>output_MAC_21_12);

	MAC_21_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_13, data_out=>output_MAC_21_13);

	MAC_21_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_14, data_out=>output_MAC_21_14);

	MAC_21_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_15, data_out=>output_MAC_21_15);

	MAC_21_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_16, data_out=>output_MAC_21_16);

	MAC_21_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_17, data_out=>output_MAC_21_17);

	MAC_21_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_18, data_out=>output_MAC_21_18);

	MAC_21_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_19, data_out=>output_MAC_21_19);

	MAC_21_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_20, data_out=>output_MAC_21_20);

	MAC_21_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_21, data_out=>output_MAC_21_21);

	MAC_21_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_22, data_out=>output_MAC_21_22);

	MAC_21_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_23, data_out=>output_MAC_21_23);

	MAC_21_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_24, data_out=>output_MAC_21_24);

	MAC_21_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_25, data_out=>output_MAC_21_25);

	MAC_21_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_26, data_out=>output_MAC_21_26);

	MAC_21_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_27, data_out=>output_MAC_21_27);

	MAC_21_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_28, data_out=>output_MAC_21_28);

	MAC_21_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_29, data_out=>output_MAC_21_29);

	MAC_21_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_30, data_out=>output_MAC_21_30);

	MAC_21_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_31, data_out=>output_MAC_21_31);

	MAC_22_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_0, data_out=>output_MAC_22_0);

	MAC_22_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_1, data_out=>output_MAC_22_1);

	MAC_22_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_2, data_out=>output_MAC_22_2);

	MAC_22_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_3, data_out=>output_MAC_22_3);

	MAC_22_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_4, data_out=>output_MAC_22_4);

	MAC_22_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_5, data_out=>output_MAC_22_5);

	MAC_22_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_6, data_out=>output_MAC_22_6);

	MAC_22_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_7, data_out=>output_MAC_22_7);

	MAC_22_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_8, data_out=>output_MAC_22_8);

	MAC_22_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_9, data_out=>output_MAC_22_9);

	MAC_22_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_10, data_out=>output_MAC_22_10);

	MAC_22_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_11, data_out=>output_MAC_22_11);

	MAC_22_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_12, data_out=>output_MAC_22_12);

	MAC_22_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_13, data_out=>output_MAC_22_13);

	MAC_22_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_14, data_out=>output_MAC_22_14);

	MAC_22_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_15, data_out=>output_MAC_22_15);

	MAC_22_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_16, data_out=>output_MAC_22_16);

	MAC_22_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_17, data_out=>output_MAC_22_17);

	MAC_22_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_18, data_out=>output_MAC_22_18);

	MAC_22_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_19, data_out=>output_MAC_22_19);

	MAC_22_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_20, data_out=>output_MAC_22_20);

	MAC_22_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_21, data_out=>output_MAC_22_21);

	MAC_22_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_22, data_out=>output_MAC_22_22);

	MAC_22_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_23, data_out=>output_MAC_22_23);

	MAC_22_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_24, data_out=>output_MAC_22_24);

	MAC_22_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_25, data_out=>output_MAC_22_25);

	MAC_22_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_26, data_out=>output_MAC_22_26);

	MAC_22_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_27, data_out=>output_MAC_22_27);

	MAC_22_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_28, data_out=>output_MAC_22_28);

	MAC_22_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_29, data_out=>output_MAC_22_29);

	MAC_22_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_30, data_out=>output_MAC_22_30);

	MAC_22_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_31, data_out=>output_MAC_22_31);

	MAC_23_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_0, data_out=>output_MAC_23_0);

	MAC_23_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_1, data_out=>output_MAC_23_1);

	MAC_23_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_2, data_out=>output_MAC_23_2);

	MAC_23_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_3, data_out=>output_MAC_23_3);

	MAC_23_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_4, data_out=>output_MAC_23_4);

	MAC_23_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_5, data_out=>output_MAC_23_5);

	MAC_23_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_6, data_out=>output_MAC_23_6);

	MAC_23_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_7, data_out=>output_MAC_23_7);

	MAC_23_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_8, data_out=>output_MAC_23_8);

	MAC_23_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_9, data_out=>output_MAC_23_9);

	MAC_23_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_10, data_out=>output_MAC_23_10);

	MAC_23_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_11, data_out=>output_MAC_23_11);

	MAC_23_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_12, data_out=>output_MAC_23_12);

	MAC_23_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_13, data_out=>output_MAC_23_13);

	MAC_23_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_14, data_out=>output_MAC_23_14);

	MAC_23_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_15, data_out=>output_MAC_23_15);

	MAC_23_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_16, data_out=>output_MAC_23_16);

	MAC_23_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_17, data_out=>output_MAC_23_17);

	MAC_23_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_18, data_out=>output_MAC_23_18);

	MAC_23_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_19, data_out=>output_MAC_23_19);

	MAC_23_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_20, data_out=>output_MAC_23_20);

	MAC_23_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_21, data_out=>output_MAC_23_21);

	MAC_23_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_22, data_out=>output_MAC_23_22);

	MAC_23_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_23, data_out=>output_MAC_23_23);

	MAC_23_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_24, data_out=>output_MAC_23_24);

	MAC_23_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_25, data_out=>output_MAC_23_25);

	MAC_23_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_26, data_out=>output_MAC_23_26);

	MAC_23_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_27, data_out=>output_MAC_23_27);

	MAC_23_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_28, data_out=>output_MAC_23_28);

	MAC_23_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_29, data_out=>output_MAC_23_29);

	MAC_23_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_30, data_out=>output_MAC_23_30);

	MAC_23_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_31, data_out=>output_MAC_23_31);

	MAC_24_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_0, data_out=>output_MAC_24_0);

	MAC_24_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_1, data_out=>output_MAC_24_1);

	MAC_24_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_2, data_out=>output_MAC_24_2);

	MAC_24_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_3, data_out=>output_MAC_24_3);

	MAC_24_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_4, data_out=>output_MAC_24_4);

	MAC_24_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_5, data_out=>output_MAC_24_5);

	MAC_24_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_6, data_out=>output_MAC_24_6);

	MAC_24_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_7, data_out=>output_MAC_24_7);

	MAC_24_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_8, data_out=>output_MAC_24_8);

	MAC_24_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_9, data_out=>output_MAC_24_9);

	MAC_24_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_10, data_out=>output_MAC_24_10);

	MAC_24_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_11, data_out=>output_MAC_24_11);

	MAC_24_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_12, data_out=>output_MAC_24_12);

	MAC_24_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_13, data_out=>output_MAC_24_13);

	MAC_24_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_14, data_out=>output_MAC_24_14);

	MAC_24_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_15, data_out=>output_MAC_24_15);

	MAC_24_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_16, data_out=>output_MAC_24_16);

	MAC_24_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_17, data_out=>output_MAC_24_17);

	MAC_24_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_18, data_out=>output_MAC_24_18);

	MAC_24_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_19, data_out=>output_MAC_24_19);

	MAC_24_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_20, data_out=>output_MAC_24_20);

	MAC_24_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_21, data_out=>output_MAC_24_21);

	MAC_24_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_22, data_out=>output_MAC_24_22);

	MAC_24_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_23, data_out=>output_MAC_24_23);

	MAC_24_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_24, data_out=>output_MAC_24_24);

	MAC_24_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_25, data_out=>output_MAC_24_25);

	MAC_24_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_26, data_out=>output_MAC_24_26);

	MAC_24_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_27, data_out=>output_MAC_24_27);

	MAC_24_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_28, data_out=>output_MAC_24_28);

	MAC_24_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_29, data_out=>output_MAC_24_29);

	MAC_24_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_30, data_out=>output_MAC_24_30);

	MAC_24_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_31, data_out=>output_MAC_24_31);

	MAC_25_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_0, data_out=>output_MAC_25_0);

	MAC_25_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_1, data_out=>output_MAC_25_1);

	MAC_25_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_2, data_out=>output_MAC_25_2);

	MAC_25_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_3, data_out=>output_MAC_25_3);

	MAC_25_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_4, data_out=>output_MAC_25_4);

	MAC_25_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_5, data_out=>output_MAC_25_5);

	MAC_25_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_6, data_out=>output_MAC_25_6);

	MAC_25_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_7, data_out=>output_MAC_25_7);

	MAC_25_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_8, data_out=>output_MAC_25_8);

	MAC_25_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_9, data_out=>output_MAC_25_9);

	MAC_25_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_10, data_out=>output_MAC_25_10);

	MAC_25_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_11, data_out=>output_MAC_25_11);

	MAC_25_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_12, data_out=>output_MAC_25_12);

	MAC_25_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_13, data_out=>output_MAC_25_13);

	MAC_25_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_14, data_out=>output_MAC_25_14);

	MAC_25_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_15, data_out=>output_MAC_25_15);

	MAC_25_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_16, data_out=>output_MAC_25_16);

	MAC_25_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_17, data_out=>output_MAC_25_17);

	MAC_25_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_18, data_out=>output_MAC_25_18);

	MAC_25_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_19, data_out=>output_MAC_25_19);

	MAC_25_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_20, data_out=>output_MAC_25_20);

	MAC_25_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_21, data_out=>output_MAC_25_21);

	MAC_25_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_22, data_out=>output_MAC_25_22);

	MAC_25_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_23, data_out=>output_MAC_25_23);

	MAC_25_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_24, data_out=>output_MAC_25_24);

	MAC_25_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_25, data_out=>output_MAC_25_25);

	MAC_25_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_26, data_out=>output_MAC_25_26);

	MAC_25_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_27, data_out=>output_MAC_25_27);

	MAC_25_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_28, data_out=>output_MAC_25_28);

	MAC_25_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_29, data_out=>output_MAC_25_29);

	MAC_25_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_30, data_out=>output_MAC_25_30);

	MAC_25_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_31, data_out=>output_MAC_25_31);

	MAC_26_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_0, data_out=>output_MAC_26_0);

	MAC_26_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_1, data_out=>output_MAC_26_1);

	MAC_26_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_2, data_out=>output_MAC_26_2);

	MAC_26_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_3, data_out=>output_MAC_26_3);

	MAC_26_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_4, data_out=>output_MAC_26_4);

	MAC_26_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_5, data_out=>output_MAC_26_5);

	MAC_26_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_6, data_out=>output_MAC_26_6);

	MAC_26_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_7, data_out=>output_MAC_26_7);

	MAC_26_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_8, data_out=>output_MAC_26_8);

	MAC_26_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_9, data_out=>output_MAC_26_9);

	MAC_26_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_10, data_out=>output_MAC_26_10);

	MAC_26_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_11, data_out=>output_MAC_26_11);

	MAC_26_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_12, data_out=>output_MAC_26_12);

	MAC_26_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_13, data_out=>output_MAC_26_13);

	MAC_26_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_14, data_out=>output_MAC_26_14);

	MAC_26_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_15, data_out=>output_MAC_26_15);

	MAC_26_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_16, data_out=>output_MAC_26_16);

	MAC_26_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_17, data_out=>output_MAC_26_17);

	MAC_26_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_18, data_out=>output_MAC_26_18);

	MAC_26_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_19, data_out=>output_MAC_26_19);

	MAC_26_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_20, data_out=>output_MAC_26_20);

	MAC_26_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_21, data_out=>output_MAC_26_21);

	MAC_26_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_22, data_out=>output_MAC_26_22);

	MAC_26_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_23, data_out=>output_MAC_26_23);

	MAC_26_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_24, data_out=>output_MAC_26_24);

	MAC_26_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_25, data_out=>output_MAC_26_25);

	MAC_26_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_26, data_out=>output_MAC_26_26);

	MAC_26_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_27, data_out=>output_MAC_26_27);

	MAC_26_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_28, data_out=>output_MAC_26_28);

	MAC_26_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_29, data_out=>output_MAC_26_29);

	MAC_26_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_30, data_out=>output_MAC_26_30);

	MAC_26_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_31, data_out=>output_MAC_26_31);

	MAC_27_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_0, data_out=>output_MAC_27_0);

	MAC_27_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_1, data_out=>output_MAC_27_1);

	MAC_27_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_2, data_out=>output_MAC_27_2);

	MAC_27_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_3, data_out=>output_MAC_27_3);

	MAC_27_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_4, data_out=>output_MAC_27_4);

	MAC_27_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_5, data_out=>output_MAC_27_5);

	MAC_27_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_6, data_out=>output_MAC_27_6);

	MAC_27_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_7, data_out=>output_MAC_27_7);

	MAC_27_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_8, data_out=>output_MAC_27_8);

	MAC_27_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_9, data_out=>output_MAC_27_9);

	MAC_27_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_10, data_out=>output_MAC_27_10);

	MAC_27_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_11, data_out=>output_MAC_27_11);

	MAC_27_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_12, data_out=>output_MAC_27_12);

	MAC_27_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_13, data_out=>output_MAC_27_13);

	MAC_27_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_14, data_out=>output_MAC_27_14);

	MAC_27_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_15, data_out=>output_MAC_27_15);

	MAC_27_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_16, data_out=>output_MAC_27_16);

	MAC_27_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_17, data_out=>output_MAC_27_17);

	MAC_27_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_18, data_out=>output_MAC_27_18);

	MAC_27_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_19, data_out=>output_MAC_27_19);

	MAC_27_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_20, data_out=>output_MAC_27_20);

	MAC_27_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_21, data_out=>output_MAC_27_21);

	MAC_27_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_22, data_out=>output_MAC_27_22);

	MAC_27_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_23, data_out=>output_MAC_27_23);

	MAC_27_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_24, data_out=>output_MAC_27_24);

	MAC_27_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_25, data_out=>output_MAC_27_25);

	MAC_27_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_26, data_out=>output_MAC_27_26);

	MAC_27_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_27, data_out=>output_MAC_27_27);

	MAC_27_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_28, data_out=>output_MAC_27_28);

	MAC_27_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_29, data_out=>output_MAC_27_29);

	MAC_27_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_30, data_out=>output_MAC_27_30);

	MAC_27_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_31, data_out=>output_MAC_27_31);

	MAC_28_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_0, data_out=>output_MAC_28_0);

	MAC_28_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_1, data_out=>output_MAC_28_1);

	MAC_28_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_2, data_out=>output_MAC_28_2);

	MAC_28_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_3, data_out=>output_MAC_28_3);

	MAC_28_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_4, data_out=>output_MAC_28_4);

	MAC_28_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_5, data_out=>output_MAC_28_5);

	MAC_28_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_6, data_out=>output_MAC_28_6);

	MAC_28_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_7, data_out=>output_MAC_28_7);

	MAC_28_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_8, data_out=>output_MAC_28_8);

	MAC_28_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_9, data_out=>output_MAC_28_9);

	MAC_28_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_10, data_out=>output_MAC_28_10);

	MAC_28_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_11, data_out=>output_MAC_28_11);

	MAC_28_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_12, data_out=>output_MAC_28_12);

	MAC_28_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_13, data_out=>output_MAC_28_13);

	MAC_28_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_14, data_out=>output_MAC_28_14);

	MAC_28_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_15, data_out=>output_MAC_28_15);

	MAC_28_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_16, data_out=>output_MAC_28_16);

	MAC_28_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_17, data_out=>output_MAC_28_17);

	MAC_28_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_18, data_out=>output_MAC_28_18);

	MAC_28_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_19, data_out=>output_MAC_28_19);

	MAC_28_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_20, data_out=>output_MAC_28_20);

	MAC_28_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_21, data_out=>output_MAC_28_21);

	MAC_28_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_22, data_out=>output_MAC_28_22);

	MAC_28_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_23, data_out=>output_MAC_28_23);

	MAC_28_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_24, data_out=>output_MAC_28_24);

	MAC_28_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_25, data_out=>output_MAC_28_25);

	MAC_28_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_26, data_out=>output_MAC_28_26);

	MAC_28_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_27, data_out=>output_MAC_28_27);

	MAC_28_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_28, data_out=>output_MAC_28_28);

	MAC_28_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_29, data_out=>output_MAC_28_29);

	MAC_28_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_30, data_out=>output_MAC_28_30);

	MAC_28_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_31, data_out=>output_MAC_28_31);

	MAC_29_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_0, data_out=>output_MAC_29_0);

	MAC_29_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_1, data_out=>output_MAC_29_1);

	MAC_29_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_2, data_out=>output_MAC_29_2);

	MAC_29_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_3, data_out=>output_MAC_29_3);

	MAC_29_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_4, data_out=>output_MAC_29_4);

	MAC_29_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_5, data_out=>output_MAC_29_5);

	MAC_29_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_6, data_out=>output_MAC_29_6);

	MAC_29_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_7, data_out=>output_MAC_29_7);

	MAC_29_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_8, data_out=>output_MAC_29_8);

	MAC_29_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_9, data_out=>output_MAC_29_9);

	MAC_29_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_10, data_out=>output_MAC_29_10);

	MAC_29_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_11, data_out=>output_MAC_29_11);

	MAC_29_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_12, data_out=>output_MAC_29_12);

	MAC_29_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_13, data_out=>output_MAC_29_13);

	MAC_29_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_14, data_out=>output_MAC_29_14);

	MAC_29_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_15, data_out=>output_MAC_29_15);

	MAC_29_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_16, data_out=>output_MAC_29_16);

	MAC_29_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_17, data_out=>output_MAC_29_17);

	MAC_29_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_18, data_out=>output_MAC_29_18);

	MAC_29_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_19, data_out=>output_MAC_29_19);

	MAC_29_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_20, data_out=>output_MAC_29_20);

	MAC_29_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_21, data_out=>output_MAC_29_21);

	MAC_29_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_22, data_out=>output_MAC_29_22);

	MAC_29_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_23, data_out=>output_MAC_29_23);

	MAC_29_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_24, data_out=>output_MAC_29_24);

	MAC_29_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_25, data_out=>output_MAC_29_25);

	MAC_29_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_26, data_out=>output_MAC_29_26);

	MAC_29_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_27, data_out=>output_MAC_29_27);

	MAC_29_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_28, data_out=>output_MAC_29_28);

	MAC_29_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_29, data_out=>output_MAC_29_29);

	MAC_29_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_30, data_out=>output_MAC_29_30);

	MAC_29_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_31, data_out=>output_MAC_29_31);

	MAC_30_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_0, data_out=>output_MAC_30_0);

	MAC_30_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_1, data_out=>output_MAC_30_1);

	MAC_30_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_2, data_out=>output_MAC_30_2);

	MAC_30_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_3, data_out=>output_MAC_30_3);

	MAC_30_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_4, data_out=>output_MAC_30_4);

	MAC_30_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_5, data_out=>output_MAC_30_5);

	MAC_30_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_6, data_out=>output_MAC_30_6);

	MAC_30_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_7, data_out=>output_MAC_30_7);

	MAC_30_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_8, data_out=>output_MAC_30_8);

	MAC_30_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_9, data_out=>output_MAC_30_9);

	MAC_30_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_10, data_out=>output_MAC_30_10);

	MAC_30_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_11, data_out=>output_MAC_30_11);

	MAC_30_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_12, data_out=>output_MAC_30_12);

	MAC_30_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_13, data_out=>output_MAC_30_13);

	MAC_30_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_14, data_out=>output_MAC_30_14);

	MAC_30_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_15, data_out=>output_MAC_30_15);

	MAC_30_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_16, data_out=>output_MAC_30_16);

	MAC_30_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_17, data_out=>output_MAC_30_17);

	MAC_30_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_18, data_out=>output_MAC_30_18);

	MAC_30_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_19, data_out=>output_MAC_30_19);

	MAC_30_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_20, data_out=>output_MAC_30_20);

	MAC_30_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_21, data_out=>output_MAC_30_21);

	MAC_30_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_22, data_out=>output_MAC_30_22);

	MAC_30_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_23, data_out=>output_MAC_30_23);

	MAC_30_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_24, data_out=>output_MAC_30_24);

	MAC_30_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_25, data_out=>output_MAC_30_25);

	MAC_30_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_26, data_out=>output_MAC_30_26);

	MAC_30_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_27, data_out=>output_MAC_30_27);

	MAC_30_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_28, data_out=>output_MAC_30_28);

	MAC_30_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_29, data_out=>output_MAC_30_29);

	MAC_30_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_30, data_out=>output_MAC_30_30);

	MAC_30_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_31, data_out=>output_MAC_30_31);

	MAC_31_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_0, data_out=>output_MAC_31_0);

	MAC_31_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_1, data_out=>output_MAC_31_1);

	MAC_31_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_2, data_out=>output_MAC_31_2);

	MAC_31_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_3, data_out=>output_MAC_31_3);

	MAC_31_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_4, data_out=>output_MAC_31_4);

	MAC_31_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_5, data_out=>output_MAC_31_5);

	MAC_31_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_6, data_out=>output_MAC_31_6);

	MAC_31_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_7, data_out=>output_MAC_31_7);

	MAC_31_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_8, data_out=>output_MAC_31_8);

	MAC_31_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_9, data_out=>output_MAC_31_9);

	MAC_31_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_10, data_out=>output_MAC_31_10);

	MAC_31_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_11, data_out=>output_MAC_31_11);

	MAC_31_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_12, data_out=>output_MAC_31_12);

	MAC_31_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_13, data_out=>output_MAC_31_13);

	MAC_31_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_14, data_out=>output_MAC_31_14);

	MAC_31_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_15, data_out=>output_MAC_31_15);

	MAC_31_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_16, data_out=>output_MAC_31_16);

	MAC_31_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_17, data_out=>output_MAC_31_17);

	MAC_31_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_18, data_out=>output_MAC_31_18);

	MAC_31_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_19, data_out=>output_MAC_31_19);

	MAC_31_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_20, data_out=>output_MAC_31_20);

	MAC_31_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_21, data_out=>output_MAC_31_21);

	MAC_31_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_22, data_out=>output_MAC_31_22);

	MAC_31_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_23, data_out=>output_MAC_31_23);

	MAC_31_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_24, data_out=>output_MAC_31_24);

	MAC_31_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_25, data_out=>output_MAC_31_25);

	MAC_31_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_26, data_out=>output_MAC_31_26);

	MAC_31_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_27, data_out=>output_MAC_31_27);

	MAC_31_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_28, data_out=>output_MAC_31_28);

	MAC_31_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_29, data_out=>output_MAC_31_29);

	MAC_31_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_30, data_out=>output_MAC_31_30);

	MAC_31_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_31, data_out=>output_MAC_31_31);

	MAC_32_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_0, data_out=>output_MAC_32_0);

	MAC_32_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_1, data_out=>output_MAC_32_1);

	MAC_32_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_2, data_out=>output_MAC_32_2);

	MAC_32_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_3, data_out=>output_MAC_32_3);

	MAC_32_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_4, data_out=>output_MAC_32_4);

	MAC_32_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_5, data_out=>output_MAC_32_5);

	MAC_32_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_6, data_out=>output_MAC_32_6);

	MAC_32_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_7, data_out=>output_MAC_32_7);

	MAC_32_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_8, data_out=>output_MAC_32_8);

	MAC_32_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_9, data_out=>output_MAC_32_9);

	MAC_32_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_10, data_out=>output_MAC_32_10);

	MAC_32_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_11, data_out=>output_MAC_32_11);

	MAC_32_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_12, data_out=>output_MAC_32_12);

	MAC_32_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_13, data_out=>output_MAC_32_13);

	MAC_32_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_14, data_out=>output_MAC_32_14);

	MAC_32_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_15, data_out=>output_MAC_32_15);

	MAC_32_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_16, data_out=>output_MAC_32_16);

	MAC_32_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_17, data_out=>output_MAC_32_17);

	MAC_32_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_18, data_out=>output_MAC_32_18);

	MAC_32_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_19, data_out=>output_MAC_32_19);

	MAC_32_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_20, data_out=>output_MAC_32_20);

	MAC_32_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_21, data_out=>output_MAC_32_21);

	MAC_32_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_22, data_out=>output_MAC_32_22);

	MAC_32_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_23, data_out=>output_MAC_32_23);

	MAC_32_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_24, data_out=>output_MAC_32_24);

	MAC_32_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_25, data_out=>output_MAC_32_25);

	MAC_32_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_26, data_out=>output_MAC_32_26);

	MAC_32_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_27, data_out=>output_MAC_32_27);

	MAC_32_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_28, data_out=>output_MAC_32_28);

	MAC_32_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_29, data_out=>output_MAC_32_29);

	MAC_32_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_30, data_out=>output_MAC_32_30);

	MAC_32_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_32, data_in_B=>reg_input_col_31, data_out=>output_MAC_32_31);

	MAC_33_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_0, data_out=>output_MAC_33_0);

	MAC_33_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_1, data_out=>output_MAC_33_1);

	MAC_33_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_2, data_out=>output_MAC_33_2);

	MAC_33_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_3, data_out=>output_MAC_33_3);

	MAC_33_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_4, data_out=>output_MAC_33_4);

	MAC_33_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_5, data_out=>output_MAC_33_5);

	MAC_33_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_6, data_out=>output_MAC_33_6);

	MAC_33_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_7, data_out=>output_MAC_33_7);

	MAC_33_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_8, data_out=>output_MAC_33_8);

	MAC_33_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_9, data_out=>output_MAC_33_9);

	MAC_33_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_10, data_out=>output_MAC_33_10);

	MAC_33_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_11, data_out=>output_MAC_33_11);

	MAC_33_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_12, data_out=>output_MAC_33_12);

	MAC_33_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_13, data_out=>output_MAC_33_13);

	MAC_33_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_14, data_out=>output_MAC_33_14);

	MAC_33_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_15, data_out=>output_MAC_33_15);

	MAC_33_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_16, data_out=>output_MAC_33_16);

	MAC_33_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_17, data_out=>output_MAC_33_17);

	MAC_33_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_18, data_out=>output_MAC_33_18);

	MAC_33_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_19, data_out=>output_MAC_33_19);

	MAC_33_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_20, data_out=>output_MAC_33_20);

	MAC_33_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_21, data_out=>output_MAC_33_21);

	MAC_33_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_22, data_out=>output_MAC_33_22);

	MAC_33_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_23, data_out=>output_MAC_33_23);

	MAC_33_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_24, data_out=>output_MAC_33_24);

	MAC_33_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_25, data_out=>output_MAC_33_25);

	MAC_33_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_26, data_out=>output_MAC_33_26);

	MAC_33_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_27, data_out=>output_MAC_33_27);

	MAC_33_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_28, data_out=>output_MAC_33_28);

	MAC_33_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_29, data_out=>output_MAC_33_29);

	MAC_33_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_30, data_out=>output_MAC_33_30);

	MAC_33_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_33, data_in_B=>reg_input_col_31, data_out=>output_MAC_33_31);

	MAC_34_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_0, data_out=>output_MAC_34_0);

	MAC_34_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_1, data_out=>output_MAC_34_1);

	MAC_34_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_2, data_out=>output_MAC_34_2);

	MAC_34_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_3, data_out=>output_MAC_34_3);

	MAC_34_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_4, data_out=>output_MAC_34_4);

	MAC_34_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_5, data_out=>output_MAC_34_5);

	MAC_34_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_6, data_out=>output_MAC_34_6);

	MAC_34_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_7, data_out=>output_MAC_34_7);

	MAC_34_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_8, data_out=>output_MAC_34_8);

	MAC_34_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_9, data_out=>output_MAC_34_9);

	MAC_34_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_10, data_out=>output_MAC_34_10);

	MAC_34_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_11, data_out=>output_MAC_34_11);

	MAC_34_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_12, data_out=>output_MAC_34_12);

	MAC_34_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_13, data_out=>output_MAC_34_13);

	MAC_34_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_14, data_out=>output_MAC_34_14);

	MAC_34_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_15, data_out=>output_MAC_34_15);

	MAC_34_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_16, data_out=>output_MAC_34_16);

	MAC_34_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_17, data_out=>output_MAC_34_17);

	MAC_34_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_18, data_out=>output_MAC_34_18);

	MAC_34_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_19, data_out=>output_MAC_34_19);

	MAC_34_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_20, data_out=>output_MAC_34_20);

	MAC_34_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_21, data_out=>output_MAC_34_21);

	MAC_34_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_22, data_out=>output_MAC_34_22);

	MAC_34_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_23, data_out=>output_MAC_34_23);

	MAC_34_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_24, data_out=>output_MAC_34_24);

	MAC_34_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_25, data_out=>output_MAC_34_25);

	MAC_34_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_26, data_out=>output_MAC_34_26);

	MAC_34_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_27, data_out=>output_MAC_34_27);

	MAC_34_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_28, data_out=>output_MAC_34_28);

	MAC_34_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_29, data_out=>output_MAC_34_29);

	MAC_34_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_30, data_out=>output_MAC_34_30);

	MAC_34_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_34, data_in_B=>reg_input_col_31, data_out=>output_MAC_34_31);

	MAC_35_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_0, data_out=>output_MAC_35_0);

	MAC_35_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_1, data_out=>output_MAC_35_1);

	MAC_35_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_2, data_out=>output_MAC_35_2);

	MAC_35_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_3, data_out=>output_MAC_35_3);

	MAC_35_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_4, data_out=>output_MAC_35_4);

	MAC_35_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_5, data_out=>output_MAC_35_5);

	MAC_35_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_6, data_out=>output_MAC_35_6);

	MAC_35_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_7, data_out=>output_MAC_35_7);

	MAC_35_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_8, data_out=>output_MAC_35_8);

	MAC_35_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_9, data_out=>output_MAC_35_9);

	MAC_35_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_10, data_out=>output_MAC_35_10);

	MAC_35_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_11, data_out=>output_MAC_35_11);

	MAC_35_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_12, data_out=>output_MAC_35_12);

	MAC_35_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_13, data_out=>output_MAC_35_13);

	MAC_35_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_14, data_out=>output_MAC_35_14);

	MAC_35_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_15, data_out=>output_MAC_35_15);

	MAC_35_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_16, data_out=>output_MAC_35_16);

	MAC_35_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_17, data_out=>output_MAC_35_17);

	MAC_35_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_18, data_out=>output_MAC_35_18);

	MAC_35_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_19, data_out=>output_MAC_35_19);

	MAC_35_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_20, data_out=>output_MAC_35_20);

	MAC_35_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_21, data_out=>output_MAC_35_21);

	MAC_35_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_22, data_out=>output_MAC_35_22);

	MAC_35_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_23, data_out=>output_MAC_35_23);

	MAC_35_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_24, data_out=>output_MAC_35_24);

	MAC_35_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_25, data_out=>output_MAC_35_25);

	MAC_35_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_26, data_out=>output_MAC_35_26);

	MAC_35_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_27, data_out=>output_MAC_35_27);

	MAC_35_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_28, data_out=>output_MAC_35_28);

	MAC_35_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_29, data_out=>output_MAC_35_29);

	MAC_35_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_30, data_out=>output_MAC_35_30);

	MAC_35_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_35, data_in_B=>reg_input_col_31, data_out=>output_MAC_35_31);

	MAC_36_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_0, data_out=>output_MAC_36_0);

	MAC_36_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_1, data_out=>output_MAC_36_1);

	MAC_36_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_2, data_out=>output_MAC_36_2);

	MAC_36_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_3, data_out=>output_MAC_36_3);

	MAC_36_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_4, data_out=>output_MAC_36_4);

	MAC_36_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_5, data_out=>output_MAC_36_5);

	MAC_36_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_6, data_out=>output_MAC_36_6);

	MAC_36_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_7, data_out=>output_MAC_36_7);

	MAC_36_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_8, data_out=>output_MAC_36_8);

	MAC_36_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_9, data_out=>output_MAC_36_9);

	MAC_36_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_10, data_out=>output_MAC_36_10);

	MAC_36_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_11, data_out=>output_MAC_36_11);

	MAC_36_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_12, data_out=>output_MAC_36_12);

	MAC_36_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_13, data_out=>output_MAC_36_13);

	MAC_36_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_14, data_out=>output_MAC_36_14);

	MAC_36_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_15, data_out=>output_MAC_36_15);

	MAC_36_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_16, data_out=>output_MAC_36_16);

	MAC_36_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_17, data_out=>output_MAC_36_17);

	MAC_36_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_18, data_out=>output_MAC_36_18);

	MAC_36_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_19, data_out=>output_MAC_36_19);

	MAC_36_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_20, data_out=>output_MAC_36_20);

	MAC_36_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_21, data_out=>output_MAC_36_21);

	MAC_36_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_22, data_out=>output_MAC_36_22);

	MAC_36_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_23, data_out=>output_MAC_36_23);

	MAC_36_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_24, data_out=>output_MAC_36_24);

	MAC_36_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_25, data_out=>output_MAC_36_25);

	MAC_36_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_26, data_out=>output_MAC_36_26);

	MAC_36_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_27, data_out=>output_MAC_36_27);

	MAC_36_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_28, data_out=>output_MAC_36_28);

	MAC_36_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_29, data_out=>output_MAC_36_29);

	MAC_36_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_30, data_out=>output_MAC_36_30);

	MAC_36_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_36, data_in_B=>reg_input_col_31, data_out=>output_MAC_36_31);

	MAC_37_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_0, data_out=>output_MAC_37_0);

	MAC_37_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_1, data_out=>output_MAC_37_1);

	MAC_37_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_2, data_out=>output_MAC_37_2);

	MAC_37_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_3, data_out=>output_MAC_37_3);

	MAC_37_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_4, data_out=>output_MAC_37_4);

	MAC_37_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_5, data_out=>output_MAC_37_5);

	MAC_37_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_6, data_out=>output_MAC_37_6);

	MAC_37_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_7, data_out=>output_MAC_37_7);

	MAC_37_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_8, data_out=>output_MAC_37_8);

	MAC_37_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_9, data_out=>output_MAC_37_9);

	MAC_37_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_10, data_out=>output_MAC_37_10);

	MAC_37_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_11, data_out=>output_MAC_37_11);

	MAC_37_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_12, data_out=>output_MAC_37_12);

	MAC_37_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_13, data_out=>output_MAC_37_13);

	MAC_37_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_14, data_out=>output_MAC_37_14);

	MAC_37_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_15, data_out=>output_MAC_37_15);

	MAC_37_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_16, data_out=>output_MAC_37_16);

	MAC_37_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_17, data_out=>output_MAC_37_17);

	MAC_37_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_18, data_out=>output_MAC_37_18);

	MAC_37_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_19, data_out=>output_MAC_37_19);

	MAC_37_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_20, data_out=>output_MAC_37_20);

	MAC_37_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_21, data_out=>output_MAC_37_21);

	MAC_37_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_22, data_out=>output_MAC_37_22);

	MAC_37_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_23, data_out=>output_MAC_37_23);

	MAC_37_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_24, data_out=>output_MAC_37_24);

	MAC_37_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_25, data_out=>output_MAC_37_25);

	MAC_37_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_26, data_out=>output_MAC_37_26);

	MAC_37_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_27, data_out=>output_MAC_37_27);

	MAC_37_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_28, data_out=>output_MAC_37_28);

	MAC_37_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_29, data_out=>output_MAC_37_29);

	MAC_37_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_30, data_out=>output_MAC_37_30);

	MAC_37_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_37, data_in_B=>reg_input_col_31, data_out=>output_MAC_37_31);

	MAC_38_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_0, data_out=>output_MAC_38_0);

	MAC_38_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_1, data_out=>output_MAC_38_1);

	MAC_38_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_2, data_out=>output_MAC_38_2);

	MAC_38_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_3, data_out=>output_MAC_38_3);

	MAC_38_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_4, data_out=>output_MAC_38_4);

	MAC_38_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_5, data_out=>output_MAC_38_5);

	MAC_38_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_6, data_out=>output_MAC_38_6);

	MAC_38_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_7, data_out=>output_MAC_38_7);

	MAC_38_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_8, data_out=>output_MAC_38_8);

	MAC_38_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_9, data_out=>output_MAC_38_9);

	MAC_38_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_10, data_out=>output_MAC_38_10);

	MAC_38_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_11, data_out=>output_MAC_38_11);

	MAC_38_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_12, data_out=>output_MAC_38_12);

	MAC_38_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_13, data_out=>output_MAC_38_13);

	MAC_38_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_14, data_out=>output_MAC_38_14);

	MAC_38_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_15, data_out=>output_MAC_38_15);

	MAC_38_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_16, data_out=>output_MAC_38_16);

	MAC_38_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_17, data_out=>output_MAC_38_17);

	MAC_38_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_18, data_out=>output_MAC_38_18);

	MAC_38_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_19, data_out=>output_MAC_38_19);

	MAC_38_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_20, data_out=>output_MAC_38_20);

	MAC_38_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_21, data_out=>output_MAC_38_21);

	MAC_38_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_22, data_out=>output_MAC_38_22);

	MAC_38_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_23, data_out=>output_MAC_38_23);

	MAC_38_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_24, data_out=>output_MAC_38_24);

	MAC_38_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_25, data_out=>output_MAC_38_25);

	MAC_38_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_26, data_out=>output_MAC_38_26);

	MAC_38_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_27, data_out=>output_MAC_38_27);

	MAC_38_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_28, data_out=>output_MAC_38_28);

	MAC_38_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_29, data_out=>output_MAC_38_29);

	MAC_38_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_30, data_out=>output_MAC_38_30);

	MAC_38_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_38, data_in_B=>reg_input_col_31, data_out=>output_MAC_38_31);

	MAC_39_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_0, data_out=>output_MAC_39_0);

	MAC_39_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_1, data_out=>output_MAC_39_1);

	MAC_39_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_2, data_out=>output_MAC_39_2);

	MAC_39_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_3, data_out=>output_MAC_39_3);

	MAC_39_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_4, data_out=>output_MAC_39_4);

	MAC_39_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_5, data_out=>output_MAC_39_5);

	MAC_39_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_6, data_out=>output_MAC_39_6);

	MAC_39_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_7, data_out=>output_MAC_39_7);

	MAC_39_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_8, data_out=>output_MAC_39_8);

	MAC_39_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_9, data_out=>output_MAC_39_9);

	MAC_39_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_10, data_out=>output_MAC_39_10);

	MAC_39_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_11, data_out=>output_MAC_39_11);

	MAC_39_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_12, data_out=>output_MAC_39_12);

	MAC_39_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_13, data_out=>output_MAC_39_13);

	MAC_39_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_14, data_out=>output_MAC_39_14);

	MAC_39_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_15, data_out=>output_MAC_39_15);

	MAC_39_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_16, data_out=>output_MAC_39_16);

	MAC_39_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_17, data_out=>output_MAC_39_17);

	MAC_39_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_18, data_out=>output_MAC_39_18);

	MAC_39_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_19, data_out=>output_MAC_39_19);

	MAC_39_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_20, data_out=>output_MAC_39_20);

	MAC_39_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_21, data_out=>output_MAC_39_21);

	MAC_39_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_22, data_out=>output_MAC_39_22);

	MAC_39_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_23, data_out=>output_MAC_39_23);

	MAC_39_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_24, data_out=>output_MAC_39_24);

	MAC_39_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_25, data_out=>output_MAC_39_25);

	MAC_39_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_26, data_out=>output_MAC_39_26);

	MAC_39_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_27, data_out=>output_MAC_39_27);

	MAC_39_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_28, data_out=>output_MAC_39_28);

	MAC_39_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_29, data_out=>output_MAC_39_29);

	MAC_39_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_30, data_out=>output_MAC_39_30);

	MAC_39_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_39, data_in_B=>reg_input_col_31, data_out=>output_MAC_39_31);

	MAC_40_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_0, data_out=>output_MAC_40_0);

	MAC_40_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_1, data_out=>output_MAC_40_1);

	MAC_40_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_2, data_out=>output_MAC_40_2);

	MAC_40_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_3, data_out=>output_MAC_40_3);

	MAC_40_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_4, data_out=>output_MAC_40_4);

	MAC_40_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_5, data_out=>output_MAC_40_5);

	MAC_40_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_6, data_out=>output_MAC_40_6);

	MAC_40_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_7, data_out=>output_MAC_40_7);

	MAC_40_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_8, data_out=>output_MAC_40_8);

	MAC_40_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_9, data_out=>output_MAC_40_9);

	MAC_40_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_10, data_out=>output_MAC_40_10);

	MAC_40_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_11, data_out=>output_MAC_40_11);

	MAC_40_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_12, data_out=>output_MAC_40_12);

	MAC_40_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_13, data_out=>output_MAC_40_13);

	MAC_40_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_14, data_out=>output_MAC_40_14);

	MAC_40_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_15, data_out=>output_MAC_40_15);

	MAC_40_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_16, data_out=>output_MAC_40_16);

	MAC_40_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_17, data_out=>output_MAC_40_17);

	MAC_40_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_18, data_out=>output_MAC_40_18);

	MAC_40_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_19, data_out=>output_MAC_40_19);

	MAC_40_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_20, data_out=>output_MAC_40_20);

	MAC_40_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_21, data_out=>output_MAC_40_21);

	MAC_40_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_22, data_out=>output_MAC_40_22);

	MAC_40_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_23, data_out=>output_MAC_40_23);

	MAC_40_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_24, data_out=>output_MAC_40_24);

	MAC_40_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_25, data_out=>output_MAC_40_25);

	MAC_40_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_26, data_out=>output_MAC_40_26);

	MAC_40_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_27, data_out=>output_MAC_40_27);

	MAC_40_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_28, data_out=>output_MAC_40_28);

	MAC_40_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_29, data_out=>output_MAC_40_29);

	MAC_40_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_30, data_out=>output_MAC_40_30);

	MAC_40_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_40, data_in_B=>reg_input_col_31, data_out=>output_MAC_40_31);

	MAC_41_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_0, data_out=>output_MAC_41_0);

	MAC_41_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_1, data_out=>output_MAC_41_1);

	MAC_41_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_2, data_out=>output_MAC_41_2);

	MAC_41_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_3, data_out=>output_MAC_41_3);

	MAC_41_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_4, data_out=>output_MAC_41_4);

	MAC_41_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_5, data_out=>output_MAC_41_5);

	MAC_41_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_6, data_out=>output_MAC_41_6);

	MAC_41_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_7, data_out=>output_MAC_41_7);

	MAC_41_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_8, data_out=>output_MAC_41_8);

	MAC_41_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_9, data_out=>output_MAC_41_9);

	MAC_41_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_10, data_out=>output_MAC_41_10);

	MAC_41_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_11, data_out=>output_MAC_41_11);

	MAC_41_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_12, data_out=>output_MAC_41_12);

	MAC_41_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_13, data_out=>output_MAC_41_13);

	MAC_41_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_14, data_out=>output_MAC_41_14);

	MAC_41_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_15, data_out=>output_MAC_41_15);

	MAC_41_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_16, data_out=>output_MAC_41_16);

	MAC_41_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_17, data_out=>output_MAC_41_17);

	MAC_41_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_18, data_out=>output_MAC_41_18);

	MAC_41_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_19, data_out=>output_MAC_41_19);

	MAC_41_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_20, data_out=>output_MAC_41_20);

	MAC_41_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_21, data_out=>output_MAC_41_21);

	MAC_41_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_22, data_out=>output_MAC_41_22);

	MAC_41_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_23, data_out=>output_MAC_41_23);

	MAC_41_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_24, data_out=>output_MAC_41_24);

	MAC_41_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_25, data_out=>output_MAC_41_25);

	MAC_41_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_26, data_out=>output_MAC_41_26);

	MAC_41_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_27, data_out=>output_MAC_41_27);

	MAC_41_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_28, data_out=>output_MAC_41_28);

	MAC_41_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_29, data_out=>output_MAC_41_29);

	MAC_41_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_30, data_out=>output_MAC_41_30);

	MAC_41_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_41, data_in_B=>reg_input_col_31, data_out=>output_MAC_41_31);

	MAC_42_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_0, data_out=>output_MAC_42_0);

	MAC_42_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_1, data_out=>output_MAC_42_1);

	MAC_42_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_2, data_out=>output_MAC_42_2);

	MAC_42_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_3, data_out=>output_MAC_42_3);

	MAC_42_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_4, data_out=>output_MAC_42_4);

	MAC_42_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_5, data_out=>output_MAC_42_5);

	MAC_42_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_6, data_out=>output_MAC_42_6);

	MAC_42_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_7, data_out=>output_MAC_42_7);

	MAC_42_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_8, data_out=>output_MAC_42_8);

	MAC_42_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_9, data_out=>output_MAC_42_9);

	MAC_42_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_10, data_out=>output_MAC_42_10);

	MAC_42_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_11, data_out=>output_MAC_42_11);

	MAC_42_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_12, data_out=>output_MAC_42_12);

	MAC_42_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_13, data_out=>output_MAC_42_13);

	MAC_42_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_14, data_out=>output_MAC_42_14);

	MAC_42_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_15, data_out=>output_MAC_42_15);

	MAC_42_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_16, data_out=>output_MAC_42_16);

	MAC_42_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_17, data_out=>output_MAC_42_17);

	MAC_42_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_18, data_out=>output_MAC_42_18);

	MAC_42_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_19, data_out=>output_MAC_42_19);

	MAC_42_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_20, data_out=>output_MAC_42_20);

	MAC_42_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_21, data_out=>output_MAC_42_21);

	MAC_42_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_22, data_out=>output_MAC_42_22);

	MAC_42_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_23, data_out=>output_MAC_42_23);

	MAC_42_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_24, data_out=>output_MAC_42_24);

	MAC_42_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_25, data_out=>output_MAC_42_25);

	MAC_42_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_26, data_out=>output_MAC_42_26);

	MAC_42_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_27, data_out=>output_MAC_42_27);

	MAC_42_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_28, data_out=>output_MAC_42_28);

	MAC_42_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_29, data_out=>output_MAC_42_29);

	MAC_42_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_30, data_out=>output_MAC_42_30);

	MAC_42_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_42, data_in_B=>reg_input_col_31, data_out=>output_MAC_42_31);

	MAC_43_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_0, data_out=>output_MAC_43_0);

	MAC_43_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_1, data_out=>output_MAC_43_1);

	MAC_43_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_2, data_out=>output_MAC_43_2);

	MAC_43_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_3, data_out=>output_MAC_43_3);

	MAC_43_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_4, data_out=>output_MAC_43_4);

	MAC_43_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_5, data_out=>output_MAC_43_5);

	MAC_43_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_6, data_out=>output_MAC_43_6);

	MAC_43_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_7, data_out=>output_MAC_43_7);

	MAC_43_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_8, data_out=>output_MAC_43_8);

	MAC_43_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_9, data_out=>output_MAC_43_9);

	MAC_43_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_10, data_out=>output_MAC_43_10);

	MAC_43_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_11, data_out=>output_MAC_43_11);

	MAC_43_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_12, data_out=>output_MAC_43_12);

	MAC_43_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_13, data_out=>output_MAC_43_13);

	MAC_43_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_14, data_out=>output_MAC_43_14);

	MAC_43_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_15, data_out=>output_MAC_43_15);

	MAC_43_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_16, data_out=>output_MAC_43_16);

	MAC_43_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_17, data_out=>output_MAC_43_17);

	MAC_43_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_18, data_out=>output_MAC_43_18);

	MAC_43_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_19, data_out=>output_MAC_43_19);

	MAC_43_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_20, data_out=>output_MAC_43_20);

	MAC_43_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_21, data_out=>output_MAC_43_21);

	MAC_43_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_22, data_out=>output_MAC_43_22);

	MAC_43_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_23, data_out=>output_MAC_43_23);

	MAC_43_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_24, data_out=>output_MAC_43_24);

	MAC_43_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_25, data_out=>output_MAC_43_25);

	MAC_43_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_26, data_out=>output_MAC_43_26);

	MAC_43_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_27, data_out=>output_MAC_43_27);

	MAC_43_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_28, data_out=>output_MAC_43_28);

	MAC_43_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_29, data_out=>output_MAC_43_29);

	MAC_43_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_30, data_out=>output_MAC_43_30);

	MAC_43_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_43, data_in_B=>reg_input_col_31, data_out=>output_MAC_43_31);

	MAC_44_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_0, data_out=>output_MAC_44_0);

	MAC_44_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_1, data_out=>output_MAC_44_1);

	MAC_44_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_2, data_out=>output_MAC_44_2);

	MAC_44_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_3, data_out=>output_MAC_44_3);

	MAC_44_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_4, data_out=>output_MAC_44_4);

	MAC_44_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_5, data_out=>output_MAC_44_5);

	MAC_44_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_6, data_out=>output_MAC_44_6);

	MAC_44_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_7, data_out=>output_MAC_44_7);

	MAC_44_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_8, data_out=>output_MAC_44_8);

	MAC_44_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_9, data_out=>output_MAC_44_9);

	MAC_44_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_10, data_out=>output_MAC_44_10);

	MAC_44_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_11, data_out=>output_MAC_44_11);

	MAC_44_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_12, data_out=>output_MAC_44_12);

	MAC_44_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_13, data_out=>output_MAC_44_13);

	MAC_44_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_14, data_out=>output_MAC_44_14);

	MAC_44_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_15, data_out=>output_MAC_44_15);

	MAC_44_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_16, data_out=>output_MAC_44_16);

	MAC_44_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_17, data_out=>output_MAC_44_17);

	MAC_44_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_18, data_out=>output_MAC_44_18);

	MAC_44_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_19, data_out=>output_MAC_44_19);

	MAC_44_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_20, data_out=>output_MAC_44_20);

	MAC_44_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_21, data_out=>output_MAC_44_21);

	MAC_44_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_22, data_out=>output_MAC_44_22);

	MAC_44_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_23, data_out=>output_MAC_44_23);

	MAC_44_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_24, data_out=>output_MAC_44_24);

	MAC_44_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_25, data_out=>output_MAC_44_25);

	MAC_44_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_26, data_out=>output_MAC_44_26);

	MAC_44_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_27, data_out=>output_MAC_44_27);

	MAC_44_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_28, data_out=>output_MAC_44_28);

	MAC_44_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_29, data_out=>output_MAC_44_29);

	MAC_44_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_30, data_out=>output_MAC_44_30);

	MAC_44_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_44, data_in_B=>reg_input_col_31, data_out=>output_MAC_44_31);

	MAC_45_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_0, data_out=>output_MAC_45_0);

	MAC_45_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_1, data_out=>output_MAC_45_1);

	MAC_45_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_2, data_out=>output_MAC_45_2);

	MAC_45_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_3, data_out=>output_MAC_45_3);

	MAC_45_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_4, data_out=>output_MAC_45_4);

	MAC_45_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_5, data_out=>output_MAC_45_5);

	MAC_45_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_6, data_out=>output_MAC_45_6);

	MAC_45_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_7, data_out=>output_MAC_45_7);

	MAC_45_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_8, data_out=>output_MAC_45_8);

	MAC_45_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_9, data_out=>output_MAC_45_9);

	MAC_45_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_10, data_out=>output_MAC_45_10);

	MAC_45_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_11, data_out=>output_MAC_45_11);

	MAC_45_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_12, data_out=>output_MAC_45_12);

	MAC_45_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_13, data_out=>output_MAC_45_13);

	MAC_45_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_14, data_out=>output_MAC_45_14);

	MAC_45_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_15, data_out=>output_MAC_45_15);

	MAC_45_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_16, data_out=>output_MAC_45_16);

	MAC_45_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_17, data_out=>output_MAC_45_17);

	MAC_45_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_18, data_out=>output_MAC_45_18);

	MAC_45_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_19, data_out=>output_MAC_45_19);

	MAC_45_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_20, data_out=>output_MAC_45_20);

	MAC_45_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_21, data_out=>output_MAC_45_21);

	MAC_45_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_22, data_out=>output_MAC_45_22);

	MAC_45_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_23, data_out=>output_MAC_45_23);

	MAC_45_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_24, data_out=>output_MAC_45_24);

	MAC_45_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_25, data_out=>output_MAC_45_25);

	MAC_45_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_26, data_out=>output_MAC_45_26);

	MAC_45_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_27, data_out=>output_MAC_45_27);

	MAC_45_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_28, data_out=>output_MAC_45_28);

	MAC_45_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_29, data_out=>output_MAC_45_29);

	MAC_45_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_30, data_out=>output_MAC_45_30);

	MAC_45_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_45, data_in_B=>reg_input_col_31, data_out=>output_MAC_45_31);

	MAC_46_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_0, data_out=>output_MAC_46_0);

	MAC_46_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_1, data_out=>output_MAC_46_1);

	MAC_46_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_2, data_out=>output_MAC_46_2);

	MAC_46_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_3, data_out=>output_MAC_46_3);

	MAC_46_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_4, data_out=>output_MAC_46_4);

	MAC_46_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_5, data_out=>output_MAC_46_5);

	MAC_46_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_6, data_out=>output_MAC_46_6);

	MAC_46_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_7, data_out=>output_MAC_46_7);

	MAC_46_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_8, data_out=>output_MAC_46_8);

	MAC_46_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_9, data_out=>output_MAC_46_9);

	MAC_46_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_10, data_out=>output_MAC_46_10);

	MAC_46_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_11, data_out=>output_MAC_46_11);

	MAC_46_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_12, data_out=>output_MAC_46_12);

	MAC_46_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_13, data_out=>output_MAC_46_13);

	MAC_46_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_14, data_out=>output_MAC_46_14);

	MAC_46_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_15, data_out=>output_MAC_46_15);

	MAC_46_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_16, data_out=>output_MAC_46_16);

	MAC_46_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_17, data_out=>output_MAC_46_17);

	MAC_46_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_18, data_out=>output_MAC_46_18);

	MAC_46_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_19, data_out=>output_MAC_46_19);

	MAC_46_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_20, data_out=>output_MAC_46_20);

	MAC_46_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_21, data_out=>output_MAC_46_21);

	MAC_46_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_22, data_out=>output_MAC_46_22);

	MAC_46_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_23, data_out=>output_MAC_46_23);

	MAC_46_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_24, data_out=>output_MAC_46_24);

	MAC_46_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_25, data_out=>output_MAC_46_25);

	MAC_46_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_26, data_out=>output_MAC_46_26);

	MAC_46_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_27, data_out=>output_MAC_46_27);

	MAC_46_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_28, data_out=>output_MAC_46_28);

	MAC_46_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_29, data_out=>output_MAC_46_29);

	MAC_46_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_30, data_out=>output_MAC_46_30);

	MAC_46_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_46, data_in_B=>reg_input_col_31, data_out=>output_MAC_46_31);

	MAC_47_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_0, data_out=>output_MAC_47_0);

	MAC_47_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_1, data_out=>output_MAC_47_1);

	MAC_47_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_2, data_out=>output_MAC_47_2);

	MAC_47_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_3, data_out=>output_MAC_47_3);

	MAC_47_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_4, data_out=>output_MAC_47_4);

	MAC_47_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_5, data_out=>output_MAC_47_5);

	MAC_47_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_6, data_out=>output_MAC_47_6);

	MAC_47_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_7, data_out=>output_MAC_47_7);

	MAC_47_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_8, data_out=>output_MAC_47_8);

	MAC_47_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_9, data_out=>output_MAC_47_9);

	MAC_47_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_10, data_out=>output_MAC_47_10);

	MAC_47_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_11, data_out=>output_MAC_47_11);

	MAC_47_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_12, data_out=>output_MAC_47_12);

	MAC_47_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_13, data_out=>output_MAC_47_13);

	MAC_47_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_14, data_out=>output_MAC_47_14);

	MAC_47_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_15, data_out=>output_MAC_47_15);

	MAC_47_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_16, data_out=>output_MAC_47_16);

	MAC_47_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_17, data_out=>output_MAC_47_17);

	MAC_47_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_18, data_out=>output_MAC_47_18);

	MAC_47_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_19, data_out=>output_MAC_47_19);

	MAC_47_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_20, data_out=>output_MAC_47_20);

	MAC_47_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_21, data_out=>output_MAC_47_21);

	MAC_47_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_22, data_out=>output_MAC_47_22);

	MAC_47_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_23, data_out=>output_MAC_47_23);

	MAC_47_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_24, data_out=>output_MAC_47_24);

	MAC_47_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_25, data_out=>output_MAC_47_25);

	MAC_47_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_26, data_out=>output_MAC_47_26);

	MAC_47_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_27, data_out=>output_MAC_47_27);

	MAC_47_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_28, data_out=>output_MAC_47_28);

	MAC_47_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_29, data_out=>output_MAC_47_29);

	MAC_47_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_30, data_out=>output_MAC_47_30);

	MAC_47_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_47, data_in_B=>reg_input_col_31, data_out=>output_MAC_47_31);

	MAC_48_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_0, data_out=>output_MAC_48_0);

	MAC_48_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_1, data_out=>output_MAC_48_1);

	MAC_48_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_2, data_out=>output_MAC_48_2);

	MAC_48_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_3, data_out=>output_MAC_48_3);

	MAC_48_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_4, data_out=>output_MAC_48_4);

	MAC_48_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_5, data_out=>output_MAC_48_5);

	MAC_48_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_6, data_out=>output_MAC_48_6);

	MAC_48_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_7, data_out=>output_MAC_48_7);

	MAC_48_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_8, data_out=>output_MAC_48_8);

	MAC_48_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_9, data_out=>output_MAC_48_9);

	MAC_48_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_10, data_out=>output_MAC_48_10);

	MAC_48_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_11, data_out=>output_MAC_48_11);

	MAC_48_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_12, data_out=>output_MAC_48_12);

	MAC_48_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_13, data_out=>output_MAC_48_13);

	MAC_48_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_14, data_out=>output_MAC_48_14);

	MAC_48_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_15, data_out=>output_MAC_48_15);

	MAC_48_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_16, data_out=>output_MAC_48_16);

	MAC_48_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_17, data_out=>output_MAC_48_17);

	MAC_48_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_18, data_out=>output_MAC_48_18);

	MAC_48_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_19, data_out=>output_MAC_48_19);

	MAC_48_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_20, data_out=>output_MAC_48_20);

	MAC_48_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_21, data_out=>output_MAC_48_21);

	MAC_48_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_22, data_out=>output_MAC_48_22);

	MAC_48_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_23, data_out=>output_MAC_48_23);

	MAC_48_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_24, data_out=>output_MAC_48_24);

	MAC_48_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_25, data_out=>output_MAC_48_25);

	MAC_48_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_26, data_out=>output_MAC_48_26);

	MAC_48_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_27, data_out=>output_MAC_48_27);

	MAC_48_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_28, data_out=>output_MAC_48_28);

	MAC_48_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_29, data_out=>output_MAC_48_29);

	MAC_48_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_30, data_out=>output_MAC_48_30);

	MAC_48_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_48, data_in_B=>reg_input_col_31, data_out=>output_MAC_48_31);

	MAC_49_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_0, data_out=>output_MAC_49_0);

	MAC_49_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_1, data_out=>output_MAC_49_1);

	MAC_49_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_2, data_out=>output_MAC_49_2);

	MAC_49_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_3, data_out=>output_MAC_49_3);

	MAC_49_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_4, data_out=>output_MAC_49_4);

	MAC_49_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_5, data_out=>output_MAC_49_5);

	MAC_49_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_6, data_out=>output_MAC_49_6);

	MAC_49_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_7, data_out=>output_MAC_49_7);

	MAC_49_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_8, data_out=>output_MAC_49_8);

	MAC_49_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_9, data_out=>output_MAC_49_9);

	MAC_49_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_10, data_out=>output_MAC_49_10);

	MAC_49_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_11, data_out=>output_MAC_49_11);

	MAC_49_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_12, data_out=>output_MAC_49_12);

	MAC_49_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_13, data_out=>output_MAC_49_13);

	MAC_49_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_14, data_out=>output_MAC_49_14);

	MAC_49_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_15, data_out=>output_MAC_49_15);

	MAC_49_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_16, data_out=>output_MAC_49_16);

	MAC_49_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_17, data_out=>output_MAC_49_17);

	MAC_49_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_18, data_out=>output_MAC_49_18);

	MAC_49_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_19, data_out=>output_MAC_49_19);

	MAC_49_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_20, data_out=>output_MAC_49_20);

	MAC_49_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_21, data_out=>output_MAC_49_21);

	MAC_49_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_22, data_out=>output_MAC_49_22);

	MAC_49_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_23, data_out=>output_MAC_49_23);

	MAC_49_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_24, data_out=>output_MAC_49_24);

	MAC_49_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_25, data_out=>output_MAC_49_25);

	MAC_49_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_26, data_out=>output_MAC_49_26);

	MAC_49_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_27, data_out=>output_MAC_49_27);

	MAC_49_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_28, data_out=>output_MAC_49_28);

	MAC_49_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_29, data_out=>output_MAC_49_29);

	MAC_49_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_30, data_out=>output_MAC_49_30);

	MAC_49_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_49, data_in_B=>reg_input_col_31, data_out=>output_MAC_49_31);

	MAC_50_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_0, data_out=>output_MAC_50_0);

	MAC_50_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_1, data_out=>output_MAC_50_1);

	MAC_50_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_2, data_out=>output_MAC_50_2);

	MAC_50_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_3, data_out=>output_MAC_50_3);

	MAC_50_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_4, data_out=>output_MAC_50_4);

	MAC_50_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_5, data_out=>output_MAC_50_5);

	MAC_50_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_6, data_out=>output_MAC_50_6);

	MAC_50_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_7, data_out=>output_MAC_50_7);

	MAC_50_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_8, data_out=>output_MAC_50_8);

	MAC_50_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_9, data_out=>output_MAC_50_9);

	MAC_50_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_10, data_out=>output_MAC_50_10);

	MAC_50_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_11, data_out=>output_MAC_50_11);

	MAC_50_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_12, data_out=>output_MAC_50_12);

	MAC_50_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_13, data_out=>output_MAC_50_13);

	MAC_50_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_14, data_out=>output_MAC_50_14);

	MAC_50_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_15, data_out=>output_MAC_50_15);

	MAC_50_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_16, data_out=>output_MAC_50_16);

	MAC_50_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_17, data_out=>output_MAC_50_17);

	MAC_50_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_18, data_out=>output_MAC_50_18);

	MAC_50_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_19, data_out=>output_MAC_50_19);

	MAC_50_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_20, data_out=>output_MAC_50_20);

	MAC_50_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_21, data_out=>output_MAC_50_21);

	MAC_50_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_22, data_out=>output_MAC_50_22);

	MAC_50_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_23, data_out=>output_MAC_50_23);

	MAC_50_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_24, data_out=>output_MAC_50_24);

	MAC_50_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_25, data_out=>output_MAC_50_25);

	MAC_50_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_26, data_out=>output_MAC_50_26);

	MAC_50_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_27, data_out=>output_MAC_50_27);

	MAC_50_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_28, data_out=>output_MAC_50_28);

	MAC_50_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_29, data_out=>output_MAC_50_29);

	MAC_50_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_30, data_out=>output_MAC_50_30);

	MAC_50_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_50, data_in_B=>reg_input_col_31, data_out=>output_MAC_50_31);

	MAC_51_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_0, data_out=>output_MAC_51_0);

	MAC_51_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_1, data_out=>output_MAC_51_1);

	MAC_51_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_2, data_out=>output_MAC_51_2);

	MAC_51_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_3, data_out=>output_MAC_51_3);

	MAC_51_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_4, data_out=>output_MAC_51_4);

	MAC_51_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_5, data_out=>output_MAC_51_5);

	MAC_51_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_6, data_out=>output_MAC_51_6);

	MAC_51_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_7, data_out=>output_MAC_51_7);

	MAC_51_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_8, data_out=>output_MAC_51_8);

	MAC_51_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_9, data_out=>output_MAC_51_9);

	MAC_51_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_10, data_out=>output_MAC_51_10);

	MAC_51_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_11, data_out=>output_MAC_51_11);

	MAC_51_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_12, data_out=>output_MAC_51_12);

	MAC_51_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_13, data_out=>output_MAC_51_13);

	MAC_51_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_14, data_out=>output_MAC_51_14);

	MAC_51_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_15, data_out=>output_MAC_51_15);

	MAC_51_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_16, data_out=>output_MAC_51_16);

	MAC_51_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_17, data_out=>output_MAC_51_17);

	MAC_51_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_18, data_out=>output_MAC_51_18);

	MAC_51_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_19, data_out=>output_MAC_51_19);

	MAC_51_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_20, data_out=>output_MAC_51_20);

	MAC_51_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_21, data_out=>output_MAC_51_21);

	MAC_51_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_22, data_out=>output_MAC_51_22);

	MAC_51_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_23, data_out=>output_MAC_51_23);

	MAC_51_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_24, data_out=>output_MAC_51_24);

	MAC_51_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_25, data_out=>output_MAC_51_25);

	MAC_51_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_26, data_out=>output_MAC_51_26);

	MAC_51_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_27, data_out=>output_MAC_51_27);

	MAC_51_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_28, data_out=>output_MAC_51_28);

	MAC_51_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_29, data_out=>output_MAC_51_29);

	MAC_51_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_30, data_out=>output_MAC_51_30);

	MAC_51_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_51, data_in_B=>reg_input_col_31, data_out=>output_MAC_51_31);

	MAC_52_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_0, data_out=>output_MAC_52_0);

	MAC_52_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_1, data_out=>output_MAC_52_1);

	MAC_52_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_2, data_out=>output_MAC_52_2);

	MAC_52_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_3, data_out=>output_MAC_52_3);

	MAC_52_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_4, data_out=>output_MAC_52_4);

	MAC_52_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_5, data_out=>output_MAC_52_5);

	MAC_52_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_6, data_out=>output_MAC_52_6);

	MAC_52_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_7, data_out=>output_MAC_52_7);

	MAC_52_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_8, data_out=>output_MAC_52_8);

	MAC_52_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_9, data_out=>output_MAC_52_9);

	MAC_52_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_10, data_out=>output_MAC_52_10);

	MAC_52_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_11, data_out=>output_MAC_52_11);

	MAC_52_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_12, data_out=>output_MAC_52_12);

	MAC_52_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_13, data_out=>output_MAC_52_13);

	MAC_52_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_14, data_out=>output_MAC_52_14);

	MAC_52_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_15, data_out=>output_MAC_52_15);

	MAC_52_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_16, data_out=>output_MAC_52_16);

	MAC_52_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_17, data_out=>output_MAC_52_17);

	MAC_52_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_18, data_out=>output_MAC_52_18);

	MAC_52_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_19, data_out=>output_MAC_52_19);

	MAC_52_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_20, data_out=>output_MAC_52_20);

	MAC_52_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_21, data_out=>output_MAC_52_21);

	MAC_52_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_22, data_out=>output_MAC_52_22);

	MAC_52_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_23, data_out=>output_MAC_52_23);

	MAC_52_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_24, data_out=>output_MAC_52_24);

	MAC_52_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_25, data_out=>output_MAC_52_25);

	MAC_52_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_26, data_out=>output_MAC_52_26);

	MAC_52_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_27, data_out=>output_MAC_52_27);

	MAC_52_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_28, data_out=>output_MAC_52_28);

	MAC_52_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_29, data_out=>output_MAC_52_29);

	MAC_52_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_30, data_out=>output_MAC_52_30);

	MAC_52_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_52, data_in_B=>reg_input_col_31, data_out=>output_MAC_52_31);

	MAC_53_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_0, data_out=>output_MAC_53_0);

	MAC_53_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_1, data_out=>output_MAC_53_1);

	MAC_53_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_2, data_out=>output_MAC_53_2);

	MAC_53_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_3, data_out=>output_MAC_53_3);

	MAC_53_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_4, data_out=>output_MAC_53_4);

	MAC_53_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_5, data_out=>output_MAC_53_5);

	MAC_53_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_6, data_out=>output_MAC_53_6);

	MAC_53_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_7, data_out=>output_MAC_53_7);

	MAC_53_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_8, data_out=>output_MAC_53_8);

	MAC_53_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_9, data_out=>output_MAC_53_9);

	MAC_53_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_10, data_out=>output_MAC_53_10);

	MAC_53_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_11, data_out=>output_MAC_53_11);

	MAC_53_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_12, data_out=>output_MAC_53_12);

	MAC_53_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_13, data_out=>output_MAC_53_13);

	MAC_53_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_14, data_out=>output_MAC_53_14);

	MAC_53_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_15, data_out=>output_MAC_53_15);

	MAC_53_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_16, data_out=>output_MAC_53_16);

	MAC_53_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_17, data_out=>output_MAC_53_17);

	MAC_53_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_18, data_out=>output_MAC_53_18);

	MAC_53_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_19, data_out=>output_MAC_53_19);

	MAC_53_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_20, data_out=>output_MAC_53_20);

	MAC_53_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_21, data_out=>output_MAC_53_21);

	MAC_53_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_22, data_out=>output_MAC_53_22);

	MAC_53_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_23, data_out=>output_MAC_53_23);

	MAC_53_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_24, data_out=>output_MAC_53_24);

	MAC_53_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_25, data_out=>output_MAC_53_25);

	MAC_53_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_26, data_out=>output_MAC_53_26);

	MAC_53_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_27, data_out=>output_MAC_53_27);

	MAC_53_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_28, data_out=>output_MAC_53_28);

	MAC_53_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_29, data_out=>output_MAC_53_29);

	MAC_53_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_30, data_out=>output_MAC_53_30);

	MAC_53_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_53, data_in_B=>reg_input_col_31, data_out=>output_MAC_53_31);

	MAC_54_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_0, data_out=>output_MAC_54_0);

	MAC_54_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_1, data_out=>output_MAC_54_1);

	MAC_54_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_2, data_out=>output_MAC_54_2);

	MAC_54_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_3, data_out=>output_MAC_54_3);

	MAC_54_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_4, data_out=>output_MAC_54_4);

	MAC_54_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_5, data_out=>output_MAC_54_5);

	MAC_54_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_6, data_out=>output_MAC_54_6);

	MAC_54_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_7, data_out=>output_MAC_54_7);

	MAC_54_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_8, data_out=>output_MAC_54_8);

	MAC_54_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_9, data_out=>output_MAC_54_9);

	MAC_54_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_10, data_out=>output_MAC_54_10);

	MAC_54_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_11, data_out=>output_MAC_54_11);

	MAC_54_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_12, data_out=>output_MAC_54_12);

	MAC_54_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_13, data_out=>output_MAC_54_13);

	MAC_54_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_14, data_out=>output_MAC_54_14);

	MAC_54_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_15, data_out=>output_MAC_54_15);

	MAC_54_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_16, data_out=>output_MAC_54_16);

	MAC_54_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_17, data_out=>output_MAC_54_17);

	MAC_54_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_18, data_out=>output_MAC_54_18);

	MAC_54_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_19, data_out=>output_MAC_54_19);

	MAC_54_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_20, data_out=>output_MAC_54_20);

	MAC_54_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_21, data_out=>output_MAC_54_21);

	MAC_54_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_22, data_out=>output_MAC_54_22);

	MAC_54_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_23, data_out=>output_MAC_54_23);

	MAC_54_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_24, data_out=>output_MAC_54_24);

	MAC_54_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_25, data_out=>output_MAC_54_25);

	MAC_54_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_26, data_out=>output_MAC_54_26);

	MAC_54_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_27, data_out=>output_MAC_54_27);

	MAC_54_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_28, data_out=>output_MAC_54_28);

	MAC_54_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_29, data_out=>output_MAC_54_29);

	MAC_54_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_30, data_out=>output_MAC_54_30);

	MAC_54_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_54, data_in_B=>reg_input_col_31, data_out=>output_MAC_54_31);

	MAC_55_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_0, data_out=>output_MAC_55_0);

	MAC_55_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_1, data_out=>output_MAC_55_1);

	MAC_55_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_2, data_out=>output_MAC_55_2);

	MAC_55_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_3, data_out=>output_MAC_55_3);

	MAC_55_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_4, data_out=>output_MAC_55_4);

	MAC_55_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_5, data_out=>output_MAC_55_5);

	MAC_55_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_6, data_out=>output_MAC_55_6);

	MAC_55_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_7, data_out=>output_MAC_55_7);

	MAC_55_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_8, data_out=>output_MAC_55_8);

	MAC_55_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_9, data_out=>output_MAC_55_9);

	MAC_55_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_10, data_out=>output_MAC_55_10);

	MAC_55_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_11, data_out=>output_MAC_55_11);

	MAC_55_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_12, data_out=>output_MAC_55_12);

	MAC_55_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_13, data_out=>output_MAC_55_13);

	MAC_55_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_14, data_out=>output_MAC_55_14);

	MAC_55_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_15, data_out=>output_MAC_55_15);

	MAC_55_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_16, data_out=>output_MAC_55_16);

	MAC_55_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_17, data_out=>output_MAC_55_17);

	MAC_55_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_18, data_out=>output_MAC_55_18);

	MAC_55_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_19, data_out=>output_MAC_55_19);

	MAC_55_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_20, data_out=>output_MAC_55_20);

	MAC_55_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_21, data_out=>output_MAC_55_21);

	MAC_55_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_22, data_out=>output_MAC_55_22);

	MAC_55_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_23, data_out=>output_MAC_55_23);

	MAC_55_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_24, data_out=>output_MAC_55_24);

	MAC_55_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_25, data_out=>output_MAC_55_25);

	MAC_55_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_26, data_out=>output_MAC_55_26);

	MAC_55_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_27, data_out=>output_MAC_55_27);

	MAC_55_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_28, data_out=>output_MAC_55_28);

	MAC_55_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_29, data_out=>output_MAC_55_29);

	MAC_55_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_30, data_out=>output_MAC_55_30);

	MAC_55_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_55, data_in_B=>reg_input_col_31, data_out=>output_MAC_55_31);

	MAC_56_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_0, data_out=>output_MAC_56_0);

	MAC_56_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_1, data_out=>output_MAC_56_1);

	MAC_56_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_2, data_out=>output_MAC_56_2);

	MAC_56_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_3, data_out=>output_MAC_56_3);

	MAC_56_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_4, data_out=>output_MAC_56_4);

	MAC_56_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_5, data_out=>output_MAC_56_5);

	MAC_56_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_6, data_out=>output_MAC_56_6);

	MAC_56_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_7, data_out=>output_MAC_56_7);

	MAC_56_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_8, data_out=>output_MAC_56_8);

	MAC_56_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_9, data_out=>output_MAC_56_9);

	MAC_56_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_10, data_out=>output_MAC_56_10);

	MAC_56_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_11, data_out=>output_MAC_56_11);

	MAC_56_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_12, data_out=>output_MAC_56_12);

	MAC_56_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_13, data_out=>output_MAC_56_13);

	MAC_56_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_14, data_out=>output_MAC_56_14);

	MAC_56_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_15, data_out=>output_MAC_56_15);

	MAC_56_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_16, data_out=>output_MAC_56_16);

	MAC_56_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_17, data_out=>output_MAC_56_17);

	MAC_56_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_18, data_out=>output_MAC_56_18);

	MAC_56_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_19, data_out=>output_MAC_56_19);

	MAC_56_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_20, data_out=>output_MAC_56_20);

	MAC_56_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_21, data_out=>output_MAC_56_21);

	MAC_56_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_22, data_out=>output_MAC_56_22);

	MAC_56_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_23, data_out=>output_MAC_56_23);

	MAC_56_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_24, data_out=>output_MAC_56_24);

	MAC_56_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_25, data_out=>output_MAC_56_25);

	MAC_56_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_26, data_out=>output_MAC_56_26);

	MAC_56_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_27, data_out=>output_MAC_56_27);

	MAC_56_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_28, data_out=>output_MAC_56_28);

	MAC_56_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_29, data_out=>output_MAC_56_29);

	MAC_56_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_30, data_out=>output_MAC_56_30);

	MAC_56_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_56, data_in_B=>reg_input_col_31, data_out=>output_MAC_56_31);

	MAC_57_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_0, data_out=>output_MAC_57_0);

	MAC_57_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_1, data_out=>output_MAC_57_1);

	MAC_57_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_2, data_out=>output_MAC_57_2);

	MAC_57_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_3, data_out=>output_MAC_57_3);

	MAC_57_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_4, data_out=>output_MAC_57_4);

	MAC_57_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_5, data_out=>output_MAC_57_5);

	MAC_57_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_6, data_out=>output_MAC_57_6);

	MAC_57_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_7, data_out=>output_MAC_57_7);

	MAC_57_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_8, data_out=>output_MAC_57_8);

	MAC_57_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_9, data_out=>output_MAC_57_9);

	MAC_57_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_10, data_out=>output_MAC_57_10);

	MAC_57_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_11, data_out=>output_MAC_57_11);

	MAC_57_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_12, data_out=>output_MAC_57_12);

	MAC_57_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_13, data_out=>output_MAC_57_13);

	MAC_57_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_14, data_out=>output_MAC_57_14);

	MAC_57_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_15, data_out=>output_MAC_57_15);

	MAC_57_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_16, data_out=>output_MAC_57_16);

	MAC_57_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_17, data_out=>output_MAC_57_17);

	MAC_57_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_18, data_out=>output_MAC_57_18);

	MAC_57_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_19, data_out=>output_MAC_57_19);

	MAC_57_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_20, data_out=>output_MAC_57_20);

	MAC_57_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_21, data_out=>output_MAC_57_21);

	MAC_57_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_22, data_out=>output_MAC_57_22);

	MAC_57_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_23, data_out=>output_MAC_57_23);

	MAC_57_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_24, data_out=>output_MAC_57_24);

	MAC_57_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_25, data_out=>output_MAC_57_25);

	MAC_57_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_26, data_out=>output_MAC_57_26);

	MAC_57_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_27, data_out=>output_MAC_57_27);

	MAC_57_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_28, data_out=>output_MAC_57_28);

	MAC_57_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_29, data_out=>output_MAC_57_29);

	MAC_57_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_30, data_out=>output_MAC_57_30);

	MAC_57_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_57, data_in_B=>reg_input_col_31, data_out=>output_MAC_57_31);

	MAC_58_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_0, data_out=>output_MAC_58_0);

	MAC_58_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_1, data_out=>output_MAC_58_1);

	MAC_58_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_2, data_out=>output_MAC_58_2);

	MAC_58_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_3, data_out=>output_MAC_58_3);

	MAC_58_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_4, data_out=>output_MAC_58_4);

	MAC_58_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_5, data_out=>output_MAC_58_5);

	MAC_58_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_6, data_out=>output_MAC_58_6);

	MAC_58_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_7, data_out=>output_MAC_58_7);

	MAC_58_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_8, data_out=>output_MAC_58_8);

	MAC_58_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_9, data_out=>output_MAC_58_9);

	MAC_58_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_10, data_out=>output_MAC_58_10);

	MAC_58_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_11, data_out=>output_MAC_58_11);

	MAC_58_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_12, data_out=>output_MAC_58_12);

	MAC_58_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_13, data_out=>output_MAC_58_13);

	MAC_58_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_14, data_out=>output_MAC_58_14);

	MAC_58_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_15, data_out=>output_MAC_58_15);

	MAC_58_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_16, data_out=>output_MAC_58_16);

	MAC_58_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_17, data_out=>output_MAC_58_17);

	MAC_58_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_18, data_out=>output_MAC_58_18);

	MAC_58_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_19, data_out=>output_MAC_58_19);

	MAC_58_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_20, data_out=>output_MAC_58_20);

	MAC_58_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_21, data_out=>output_MAC_58_21);

	MAC_58_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_22, data_out=>output_MAC_58_22);

	MAC_58_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_23, data_out=>output_MAC_58_23);

	MAC_58_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_24, data_out=>output_MAC_58_24);

	MAC_58_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_25, data_out=>output_MAC_58_25);

	MAC_58_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_26, data_out=>output_MAC_58_26);

	MAC_58_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_27, data_out=>output_MAC_58_27);

	MAC_58_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_28, data_out=>output_MAC_58_28);

	MAC_58_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_29, data_out=>output_MAC_58_29);

	MAC_58_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_30, data_out=>output_MAC_58_30);

	MAC_58_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_58, data_in_B=>reg_input_col_31, data_out=>output_MAC_58_31);

	MAC_59_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_0, data_out=>output_MAC_59_0);

	MAC_59_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_1, data_out=>output_MAC_59_1);

	MAC_59_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_2, data_out=>output_MAC_59_2);

	MAC_59_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_3, data_out=>output_MAC_59_3);

	MAC_59_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_4, data_out=>output_MAC_59_4);

	MAC_59_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_5, data_out=>output_MAC_59_5);

	MAC_59_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_6, data_out=>output_MAC_59_6);

	MAC_59_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_7, data_out=>output_MAC_59_7);

	MAC_59_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_8, data_out=>output_MAC_59_8);

	MAC_59_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_9, data_out=>output_MAC_59_9);

	MAC_59_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_10, data_out=>output_MAC_59_10);

	MAC_59_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_11, data_out=>output_MAC_59_11);

	MAC_59_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_12, data_out=>output_MAC_59_12);

	MAC_59_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_13, data_out=>output_MAC_59_13);

	MAC_59_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_14, data_out=>output_MAC_59_14);

	MAC_59_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_15, data_out=>output_MAC_59_15);

	MAC_59_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_16, data_out=>output_MAC_59_16);

	MAC_59_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_17, data_out=>output_MAC_59_17);

	MAC_59_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_18, data_out=>output_MAC_59_18);

	MAC_59_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_19, data_out=>output_MAC_59_19);

	MAC_59_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_20, data_out=>output_MAC_59_20);

	MAC_59_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_21, data_out=>output_MAC_59_21);

	MAC_59_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_22, data_out=>output_MAC_59_22);

	MAC_59_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_23, data_out=>output_MAC_59_23);

	MAC_59_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_24, data_out=>output_MAC_59_24);

	MAC_59_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_25, data_out=>output_MAC_59_25);

	MAC_59_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_26, data_out=>output_MAC_59_26);

	MAC_59_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_27, data_out=>output_MAC_59_27);

	MAC_59_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_28, data_out=>output_MAC_59_28);

	MAC_59_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_29, data_out=>output_MAC_59_29);

	MAC_59_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_30, data_out=>output_MAC_59_30);

	MAC_59_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_59, data_in_B=>reg_input_col_31, data_out=>output_MAC_59_31);

	MAC_60_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_0, data_out=>output_MAC_60_0);

	MAC_60_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_1, data_out=>output_MAC_60_1);

	MAC_60_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_2, data_out=>output_MAC_60_2);

	MAC_60_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_3, data_out=>output_MAC_60_3);

	MAC_60_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_4, data_out=>output_MAC_60_4);

	MAC_60_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_5, data_out=>output_MAC_60_5);

	MAC_60_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_6, data_out=>output_MAC_60_6);

	MAC_60_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_7, data_out=>output_MAC_60_7);

	MAC_60_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_8, data_out=>output_MAC_60_8);

	MAC_60_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_9, data_out=>output_MAC_60_9);

	MAC_60_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_10, data_out=>output_MAC_60_10);

	MAC_60_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_11, data_out=>output_MAC_60_11);

	MAC_60_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_12, data_out=>output_MAC_60_12);

	MAC_60_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_13, data_out=>output_MAC_60_13);

	MAC_60_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_14, data_out=>output_MAC_60_14);

	MAC_60_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_15, data_out=>output_MAC_60_15);

	MAC_60_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_16, data_out=>output_MAC_60_16);

	MAC_60_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_17, data_out=>output_MAC_60_17);

	MAC_60_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_18, data_out=>output_MAC_60_18);

	MAC_60_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_19, data_out=>output_MAC_60_19);

	MAC_60_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_20, data_out=>output_MAC_60_20);

	MAC_60_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_21, data_out=>output_MAC_60_21);

	MAC_60_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_22, data_out=>output_MAC_60_22);

	MAC_60_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_23, data_out=>output_MAC_60_23);

	MAC_60_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_24, data_out=>output_MAC_60_24);

	MAC_60_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_25, data_out=>output_MAC_60_25);

	MAC_60_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_26, data_out=>output_MAC_60_26);

	MAC_60_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_27, data_out=>output_MAC_60_27);

	MAC_60_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_28, data_out=>output_MAC_60_28);

	MAC_60_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_29, data_out=>output_MAC_60_29);

	MAC_60_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_30, data_out=>output_MAC_60_30);

	MAC_60_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_60, data_in_B=>reg_input_col_31, data_out=>output_MAC_60_31);

	MAC_61_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_0, data_out=>output_MAC_61_0);

	MAC_61_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_1, data_out=>output_MAC_61_1);

	MAC_61_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_2, data_out=>output_MAC_61_2);

	MAC_61_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_3, data_out=>output_MAC_61_3);

	MAC_61_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_4, data_out=>output_MAC_61_4);

	MAC_61_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_5, data_out=>output_MAC_61_5);

	MAC_61_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_6, data_out=>output_MAC_61_6);

	MAC_61_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_7, data_out=>output_MAC_61_7);

	MAC_61_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_8, data_out=>output_MAC_61_8);

	MAC_61_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_9, data_out=>output_MAC_61_9);

	MAC_61_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_10, data_out=>output_MAC_61_10);

	MAC_61_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_11, data_out=>output_MAC_61_11);

	MAC_61_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_12, data_out=>output_MAC_61_12);

	MAC_61_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_13, data_out=>output_MAC_61_13);

	MAC_61_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_14, data_out=>output_MAC_61_14);

	MAC_61_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_15, data_out=>output_MAC_61_15);

	MAC_61_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_16, data_out=>output_MAC_61_16);

	MAC_61_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_17, data_out=>output_MAC_61_17);

	MAC_61_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_18, data_out=>output_MAC_61_18);

	MAC_61_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_19, data_out=>output_MAC_61_19);

	MAC_61_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_20, data_out=>output_MAC_61_20);

	MAC_61_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_21, data_out=>output_MAC_61_21);

	MAC_61_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_22, data_out=>output_MAC_61_22);

	MAC_61_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_23, data_out=>output_MAC_61_23);

	MAC_61_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_24, data_out=>output_MAC_61_24);

	MAC_61_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_25, data_out=>output_MAC_61_25);

	MAC_61_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_26, data_out=>output_MAC_61_26);

	MAC_61_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_27, data_out=>output_MAC_61_27);

	MAC_61_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_28, data_out=>output_MAC_61_28);

	MAC_61_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_29, data_out=>output_MAC_61_29);

	MAC_61_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_30, data_out=>output_MAC_61_30);

	MAC_61_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_61, data_in_B=>reg_input_col_31, data_out=>output_MAC_61_31);

	MAC_62_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_0, data_out=>output_MAC_62_0);

	MAC_62_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_1, data_out=>output_MAC_62_1);

	MAC_62_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_2, data_out=>output_MAC_62_2);

	MAC_62_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_3, data_out=>output_MAC_62_3);

	MAC_62_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_4, data_out=>output_MAC_62_4);

	MAC_62_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_5, data_out=>output_MAC_62_5);

	MAC_62_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_6, data_out=>output_MAC_62_6);

	MAC_62_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_7, data_out=>output_MAC_62_7);

	MAC_62_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_8, data_out=>output_MAC_62_8);

	MAC_62_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_9, data_out=>output_MAC_62_9);

	MAC_62_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_10, data_out=>output_MAC_62_10);

	MAC_62_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_11, data_out=>output_MAC_62_11);

	MAC_62_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_12, data_out=>output_MAC_62_12);

	MAC_62_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_13, data_out=>output_MAC_62_13);

	MAC_62_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_14, data_out=>output_MAC_62_14);

	MAC_62_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_15, data_out=>output_MAC_62_15);

	MAC_62_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_16, data_out=>output_MAC_62_16);

	MAC_62_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_17, data_out=>output_MAC_62_17);

	MAC_62_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_18, data_out=>output_MAC_62_18);

	MAC_62_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_19, data_out=>output_MAC_62_19);

	MAC_62_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_20, data_out=>output_MAC_62_20);

	MAC_62_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_21, data_out=>output_MAC_62_21);

	MAC_62_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_22, data_out=>output_MAC_62_22);

	MAC_62_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_23, data_out=>output_MAC_62_23);

	MAC_62_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_24, data_out=>output_MAC_62_24);

	MAC_62_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_25, data_out=>output_MAC_62_25);

	MAC_62_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_26, data_out=>output_MAC_62_26);

	MAC_62_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_27, data_out=>output_MAC_62_27);

	MAC_62_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_28, data_out=>output_MAC_62_28);

	MAC_62_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_29, data_out=>output_MAC_62_29);

	MAC_62_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_30, data_out=>output_MAC_62_30);

	MAC_62_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_62, data_in_B=>reg_input_col_31, data_out=>output_MAC_62_31);

	MAC_63_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_0, data_out=>output_MAC_63_0);

	MAC_63_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_1, data_out=>output_MAC_63_1);

	MAC_63_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_2, data_out=>output_MAC_63_2);

	MAC_63_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_3, data_out=>output_MAC_63_3);

	MAC_63_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_4, data_out=>output_MAC_63_4);

	MAC_63_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_5, data_out=>output_MAC_63_5);

	MAC_63_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_6, data_out=>output_MAC_63_6);

	MAC_63_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_7, data_out=>output_MAC_63_7);

	MAC_63_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_8, data_out=>output_MAC_63_8);

	MAC_63_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_9, data_out=>output_MAC_63_9);

	MAC_63_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_10, data_out=>output_MAC_63_10);

	MAC_63_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_11, data_out=>output_MAC_63_11);

	MAC_63_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_12, data_out=>output_MAC_63_12);

	MAC_63_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_13, data_out=>output_MAC_63_13);

	MAC_63_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_14, data_out=>output_MAC_63_14);

	MAC_63_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_15, data_out=>output_MAC_63_15);

	MAC_63_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_16, data_out=>output_MAC_63_16);

	MAC_63_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_17, data_out=>output_MAC_63_17);

	MAC_63_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_18, data_out=>output_MAC_63_18);

	MAC_63_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_19, data_out=>output_MAC_63_19);

	MAC_63_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_20, data_out=>output_MAC_63_20);

	MAC_63_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_21, data_out=>output_MAC_63_21);

	MAC_63_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_22, data_out=>output_MAC_63_22);

	MAC_63_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_23, data_out=>output_MAC_63_23);

	MAC_63_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_24, data_out=>output_MAC_63_24);

	MAC_63_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_25, data_out=>output_MAC_63_25);

	MAC_63_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_26, data_out=>output_MAC_63_26);

	MAC_63_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_27, data_out=>output_MAC_63_27);

	MAC_63_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_28, data_out=>output_MAC_63_28);

	MAC_63_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_29, data_out=>output_MAC_63_29);

	MAC_63_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_30, data_out=>output_MAC_63_30);

	MAC_63_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_63, data_in_B=>reg_input_col_31, data_out=>output_MAC_63_31);

	MAC_64_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_0, data_out=>output_MAC_64_0);

	MAC_64_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_1, data_out=>output_MAC_64_1);

	MAC_64_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_2, data_out=>output_MAC_64_2);

	MAC_64_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_3, data_out=>output_MAC_64_3);

	MAC_64_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_4, data_out=>output_MAC_64_4);

	MAC_64_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_5, data_out=>output_MAC_64_5);

	MAC_64_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_6, data_out=>output_MAC_64_6);

	MAC_64_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_7, data_out=>output_MAC_64_7);

	MAC_64_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_8, data_out=>output_MAC_64_8);

	MAC_64_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_9, data_out=>output_MAC_64_9);

	MAC_64_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_10, data_out=>output_MAC_64_10);

	MAC_64_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_11, data_out=>output_MAC_64_11);

	MAC_64_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_12, data_out=>output_MAC_64_12);

	MAC_64_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_13, data_out=>output_MAC_64_13);

	MAC_64_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_14, data_out=>output_MAC_64_14);

	MAC_64_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_15, data_out=>output_MAC_64_15);

	MAC_64_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_16, data_out=>output_MAC_64_16);

	MAC_64_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_17, data_out=>output_MAC_64_17);

	MAC_64_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_18, data_out=>output_MAC_64_18);

	MAC_64_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_19, data_out=>output_MAC_64_19);

	MAC_64_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_20, data_out=>output_MAC_64_20);

	MAC_64_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_21, data_out=>output_MAC_64_21);

	MAC_64_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_22, data_out=>output_MAC_64_22);

	MAC_64_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_23, data_out=>output_MAC_64_23);

	MAC_64_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_24, data_out=>output_MAC_64_24);

	MAC_64_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_25, data_out=>output_MAC_64_25);

	MAC_64_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_26, data_out=>output_MAC_64_26);

	MAC_64_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_27, data_out=>output_MAC_64_27);

	MAC_64_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_28, data_out=>output_MAC_64_28);

	MAC_64_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_29, data_out=>output_MAC_64_29);

	MAC_64_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_30, data_out=>output_MAC_64_30);

	MAC_64_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_64, data_in_B=>reg_input_col_31, data_out=>output_MAC_64_31);

	MAC_65_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_0, data_out=>output_MAC_65_0);

	MAC_65_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_1, data_out=>output_MAC_65_1);

	MAC_65_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_2, data_out=>output_MAC_65_2);

	MAC_65_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_3, data_out=>output_MAC_65_3);

	MAC_65_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_4, data_out=>output_MAC_65_4);

	MAC_65_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_5, data_out=>output_MAC_65_5);

	MAC_65_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_6, data_out=>output_MAC_65_6);

	MAC_65_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_7, data_out=>output_MAC_65_7);

	MAC_65_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_8, data_out=>output_MAC_65_8);

	MAC_65_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_9, data_out=>output_MAC_65_9);

	MAC_65_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_10, data_out=>output_MAC_65_10);

	MAC_65_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_11, data_out=>output_MAC_65_11);

	MAC_65_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_12, data_out=>output_MAC_65_12);

	MAC_65_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_13, data_out=>output_MAC_65_13);

	MAC_65_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_14, data_out=>output_MAC_65_14);

	MAC_65_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_15, data_out=>output_MAC_65_15);

	MAC_65_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_16, data_out=>output_MAC_65_16);

	MAC_65_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_17, data_out=>output_MAC_65_17);

	MAC_65_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_18, data_out=>output_MAC_65_18);

	MAC_65_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_19, data_out=>output_MAC_65_19);

	MAC_65_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_20, data_out=>output_MAC_65_20);

	MAC_65_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_21, data_out=>output_MAC_65_21);

	MAC_65_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_22, data_out=>output_MAC_65_22);

	MAC_65_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_23, data_out=>output_MAC_65_23);

	MAC_65_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_24, data_out=>output_MAC_65_24);

	MAC_65_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_25, data_out=>output_MAC_65_25);

	MAC_65_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_26, data_out=>output_MAC_65_26);

	MAC_65_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_27, data_out=>output_MAC_65_27);

	MAC_65_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_28, data_out=>output_MAC_65_28);

	MAC_65_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_29, data_out=>output_MAC_65_29);

	MAC_65_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_30, data_out=>output_MAC_65_30);

	MAC_65_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_65, data_in_B=>reg_input_col_31, data_out=>output_MAC_65_31);

	MAC_66_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_0, data_out=>output_MAC_66_0);

	MAC_66_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_1, data_out=>output_MAC_66_1);

	MAC_66_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_2, data_out=>output_MAC_66_2);

	MAC_66_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_3, data_out=>output_MAC_66_3);

	MAC_66_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_4, data_out=>output_MAC_66_4);

	MAC_66_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_5, data_out=>output_MAC_66_5);

	MAC_66_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_6, data_out=>output_MAC_66_6);

	MAC_66_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_7, data_out=>output_MAC_66_7);

	MAC_66_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_8, data_out=>output_MAC_66_8);

	MAC_66_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_9, data_out=>output_MAC_66_9);

	MAC_66_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_10, data_out=>output_MAC_66_10);

	MAC_66_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_11, data_out=>output_MAC_66_11);

	MAC_66_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_12, data_out=>output_MAC_66_12);

	MAC_66_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_13, data_out=>output_MAC_66_13);

	MAC_66_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_14, data_out=>output_MAC_66_14);

	MAC_66_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_15, data_out=>output_MAC_66_15);

	MAC_66_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_16, data_out=>output_MAC_66_16);

	MAC_66_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_17, data_out=>output_MAC_66_17);

	MAC_66_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_18, data_out=>output_MAC_66_18);

	MAC_66_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_19, data_out=>output_MAC_66_19);

	MAC_66_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_20, data_out=>output_MAC_66_20);

	MAC_66_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_21, data_out=>output_MAC_66_21);

	MAC_66_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_22, data_out=>output_MAC_66_22);

	MAC_66_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_23, data_out=>output_MAC_66_23);

	MAC_66_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_24, data_out=>output_MAC_66_24);

	MAC_66_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_25, data_out=>output_MAC_66_25);

	MAC_66_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_26, data_out=>output_MAC_66_26);

	MAC_66_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_27, data_out=>output_MAC_66_27);

	MAC_66_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_28, data_out=>output_MAC_66_28);

	MAC_66_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_29, data_out=>output_MAC_66_29);

	MAC_66_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_30, data_out=>output_MAC_66_30);

	MAC_66_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_66, data_in_B=>reg_input_col_31, data_out=>output_MAC_66_31);

	MAC_67_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_0, data_out=>output_MAC_67_0);

	MAC_67_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_1, data_out=>output_MAC_67_1);

	MAC_67_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_2, data_out=>output_MAC_67_2);

	MAC_67_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_3, data_out=>output_MAC_67_3);

	MAC_67_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_4, data_out=>output_MAC_67_4);

	MAC_67_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_5, data_out=>output_MAC_67_5);

	MAC_67_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_6, data_out=>output_MAC_67_6);

	MAC_67_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_7, data_out=>output_MAC_67_7);

	MAC_67_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_8, data_out=>output_MAC_67_8);

	MAC_67_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_9, data_out=>output_MAC_67_9);

	MAC_67_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_10, data_out=>output_MAC_67_10);

	MAC_67_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_11, data_out=>output_MAC_67_11);

	MAC_67_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_12, data_out=>output_MAC_67_12);

	MAC_67_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_13, data_out=>output_MAC_67_13);

	MAC_67_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_14, data_out=>output_MAC_67_14);

	MAC_67_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_15, data_out=>output_MAC_67_15);

	MAC_67_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_16, data_out=>output_MAC_67_16);

	MAC_67_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_17, data_out=>output_MAC_67_17);

	MAC_67_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_18, data_out=>output_MAC_67_18);

	MAC_67_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_19, data_out=>output_MAC_67_19);

	MAC_67_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_20, data_out=>output_MAC_67_20);

	MAC_67_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_21, data_out=>output_MAC_67_21);

	MAC_67_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_22, data_out=>output_MAC_67_22);

	MAC_67_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_23, data_out=>output_MAC_67_23);

	MAC_67_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_24, data_out=>output_MAC_67_24);

	MAC_67_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_25, data_out=>output_MAC_67_25);

	MAC_67_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_26, data_out=>output_MAC_67_26);

	MAC_67_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_27, data_out=>output_MAC_67_27);

	MAC_67_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_28, data_out=>output_MAC_67_28);

	MAC_67_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_29, data_out=>output_MAC_67_29);

	MAC_67_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_30, data_out=>output_MAC_67_30);

	MAC_67_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_67, data_in_B=>reg_input_col_31, data_out=>output_MAC_67_31);

	MAC_68_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_0, data_out=>output_MAC_68_0);

	MAC_68_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_1, data_out=>output_MAC_68_1);

	MAC_68_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_2, data_out=>output_MAC_68_2);

	MAC_68_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_3, data_out=>output_MAC_68_3);

	MAC_68_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_4, data_out=>output_MAC_68_4);

	MAC_68_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_5, data_out=>output_MAC_68_5);

	MAC_68_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_6, data_out=>output_MAC_68_6);

	MAC_68_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_7, data_out=>output_MAC_68_7);

	MAC_68_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_8, data_out=>output_MAC_68_8);

	MAC_68_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_9, data_out=>output_MAC_68_9);

	MAC_68_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_10, data_out=>output_MAC_68_10);

	MAC_68_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_11, data_out=>output_MAC_68_11);

	MAC_68_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_12, data_out=>output_MAC_68_12);

	MAC_68_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_13, data_out=>output_MAC_68_13);

	MAC_68_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_14, data_out=>output_MAC_68_14);

	MAC_68_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_15, data_out=>output_MAC_68_15);

	MAC_68_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_16, data_out=>output_MAC_68_16);

	MAC_68_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_17, data_out=>output_MAC_68_17);

	MAC_68_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_18, data_out=>output_MAC_68_18);

	MAC_68_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_19, data_out=>output_MAC_68_19);

	MAC_68_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_20, data_out=>output_MAC_68_20);

	MAC_68_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_21, data_out=>output_MAC_68_21);

	MAC_68_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_22, data_out=>output_MAC_68_22);

	MAC_68_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_23, data_out=>output_MAC_68_23);

	MAC_68_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_24, data_out=>output_MAC_68_24);

	MAC_68_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_25, data_out=>output_MAC_68_25);

	MAC_68_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_26, data_out=>output_MAC_68_26);

	MAC_68_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_27, data_out=>output_MAC_68_27);

	MAC_68_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_28, data_out=>output_MAC_68_28);

	MAC_68_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_29, data_out=>output_MAC_68_29);

	MAC_68_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_30, data_out=>output_MAC_68_30);

	MAC_68_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_68, data_in_B=>reg_input_col_31, data_out=>output_MAC_68_31);

	MAC_69_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_0, data_out=>output_MAC_69_0);

	MAC_69_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_1, data_out=>output_MAC_69_1);

	MAC_69_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_2, data_out=>output_MAC_69_2);

	MAC_69_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_3, data_out=>output_MAC_69_3);

	MAC_69_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_4, data_out=>output_MAC_69_4);

	MAC_69_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_5, data_out=>output_MAC_69_5);

	MAC_69_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_6, data_out=>output_MAC_69_6);

	MAC_69_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_7, data_out=>output_MAC_69_7);

	MAC_69_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_8, data_out=>output_MAC_69_8);

	MAC_69_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_9, data_out=>output_MAC_69_9);

	MAC_69_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_10, data_out=>output_MAC_69_10);

	MAC_69_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_11, data_out=>output_MAC_69_11);

	MAC_69_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_12, data_out=>output_MAC_69_12);

	MAC_69_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_13, data_out=>output_MAC_69_13);

	MAC_69_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_14, data_out=>output_MAC_69_14);

	MAC_69_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_15, data_out=>output_MAC_69_15);

	MAC_69_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_16, data_out=>output_MAC_69_16);

	MAC_69_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_17, data_out=>output_MAC_69_17);

	MAC_69_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_18, data_out=>output_MAC_69_18);

	MAC_69_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_19, data_out=>output_MAC_69_19);

	MAC_69_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_20, data_out=>output_MAC_69_20);

	MAC_69_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_21, data_out=>output_MAC_69_21);

	MAC_69_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_22, data_out=>output_MAC_69_22);

	MAC_69_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_23, data_out=>output_MAC_69_23);

	MAC_69_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_24, data_out=>output_MAC_69_24);

	MAC_69_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_25, data_out=>output_MAC_69_25);

	MAC_69_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_26, data_out=>output_MAC_69_26);

	MAC_69_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_27, data_out=>output_MAC_69_27);

	MAC_69_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_28, data_out=>output_MAC_69_28);

	MAC_69_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_29, data_out=>output_MAC_69_29);

	MAC_69_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_30, data_out=>output_MAC_69_30);

	MAC_69_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_69, data_in_B=>reg_input_col_31, data_out=>output_MAC_69_31);

	MAC_70_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_0, data_out=>output_MAC_70_0);

	MAC_70_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_1, data_out=>output_MAC_70_1);

	MAC_70_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_2, data_out=>output_MAC_70_2);

	MAC_70_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_3, data_out=>output_MAC_70_3);

	MAC_70_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_4, data_out=>output_MAC_70_4);

	MAC_70_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_5, data_out=>output_MAC_70_5);

	MAC_70_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_6, data_out=>output_MAC_70_6);

	MAC_70_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_7, data_out=>output_MAC_70_7);

	MAC_70_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_8, data_out=>output_MAC_70_8);

	MAC_70_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_9, data_out=>output_MAC_70_9);

	MAC_70_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_10, data_out=>output_MAC_70_10);

	MAC_70_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_11, data_out=>output_MAC_70_11);

	MAC_70_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_12, data_out=>output_MAC_70_12);

	MAC_70_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_13, data_out=>output_MAC_70_13);

	MAC_70_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_14, data_out=>output_MAC_70_14);

	MAC_70_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_15, data_out=>output_MAC_70_15);

	MAC_70_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_16, data_out=>output_MAC_70_16);

	MAC_70_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_17, data_out=>output_MAC_70_17);

	MAC_70_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_18, data_out=>output_MAC_70_18);

	MAC_70_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_19, data_out=>output_MAC_70_19);

	MAC_70_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_20, data_out=>output_MAC_70_20);

	MAC_70_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_21, data_out=>output_MAC_70_21);

	MAC_70_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_22, data_out=>output_MAC_70_22);

	MAC_70_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_23, data_out=>output_MAC_70_23);

	MAC_70_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_24, data_out=>output_MAC_70_24);

	MAC_70_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_25, data_out=>output_MAC_70_25);

	MAC_70_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_26, data_out=>output_MAC_70_26);

	MAC_70_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_27, data_out=>output_MAC_70_27);

	MAC_70_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_28, data_out=>output_MAC_70_28);

	MAC_70_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_29, data_out=>output_MAC_70_29);

	MAC_70_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_30, data_out=>output_MAC_70_30);

	MAC_70_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_70, data_in_B=>reg_input_col_31, data_out=>output_MAC_70_31);

	MAC_71_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_0, data_out=>output_MAC_71_0);

	MAC_71_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_1, data_out=>output_MAC_71_1);

	MAC_71_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_2, data_out=>output_MAC_71_2);

	MAC_71_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_3, data_out=>output_MAC_71_3);

	MAC_71_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_4, data_out=>output_MAC_71_4);

	MAC_71_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_5, data_out=>output_MAC_71_5);

	MAC_71_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_6, data_out=>output_MAC_71_6);

	MAC_71_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_7, data_out=>output_MAC_71_7);

	MAC_71_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_8, data_out=>output_MAC_71_8);

	MAC_71_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_9, data_out=>output_MAC_71_9);

	MAC_71_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_10, data_out=>output_MAC_71_10);

	MAC_71_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_11, data_out=>output_MAC_71_11);

	MAC_71_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_12, data_out=>output_MAC_71_12);

	MAC_71_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_13, data_out=>output_MAC_71_13);

	MAC_71_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_14, data_out=>output_MAC_71_14);

	MAC_71_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_15, data_out=>output_MAC_71_15);

	MAC_71_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_16, data_out=>output_MAC_71_16);

	MAC_71_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_17, data_out=>output_MAC_71_17);

	MAC_71_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_18, data_out=>output_MAC_71_18);

	MAC_71_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_19, data_out=>output_MAC_71_19);

	MAC_71_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_20, data_out=>output_MAC_71_20);

	MAC_71_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_21, data_out=>output_MAC_71_21);

	MAC_71_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_22, data_out=>output_MAC_71_22);

	MAC_71_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_23, data_out=>output_MAC_71_23);

	MAC_71_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_24, data_out=>output_MAC_71_24);

	MAC_71_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_25, data_out=>output_MAC_71_25);

	MAC_71_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_26, data_out=>output_MAC_71_26);

	MAC_71_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_27, data_out=>output_MAC_71_27);

	MAC_71_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_28, data_out=>output_MAC_71_28);

	MAC_71_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_29, data_out=>output_MAC_71_29);

	MAC_71_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_30, data_out=>output_MAC_71_30);

	MAC_71_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_71, data_in_B=>reg_input_col_31, data_out=>output_MAC_71_31);

	MAC_72_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_0, data_out=>output_MAC_72_0);

	MAC_72_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_1, data_out=>output_MAC_72_1);

	MAC_72_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_2, data_out=>output_MAC_72_2);

	MAC_72_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_3, data_out=>output_MAC_72_3);

	MAC_72_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_4, data_out=>output_MAC_72_4);

	MAC_72_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_5, data_out=>output_MAC_72_5);

	MAC_72_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_6, data_out=>output_MAC_72_6);

	MAC_72_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_7, data_out=>output_MAC_72_7);

	MAC_72_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_8, data_out=>output_MAC_72_8);

	MAC_72_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_9, data_out=>output_MAC_72_9);

	MAC_72_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_10, data_out=>output_MAC_72_10);

	MAC_72_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_11, data_out=>output_MAC_72_11);

	MAC_72_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_12, data_out=>output_MAC_72_12);

	MAC_72_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_13, data_out=>output_MAC_72_13);

	MAC_72_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_14, data_out=>output_MAC_72_14);

	MAC_72_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_15, data_out=>output_MAC_72_15);

	MAC_72_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_16, data_out=>output_MAC_72_16);

	MAC_72_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_17, data_out=>output_MAC_72_17);

	MAC_72_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_18, data_out=>output_MAC_72_18);

	MAC_72_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_19, data_out=>output_MAC_72_19);

	MAC_72_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_20, data_out=>output_MAC_72_20);

	MAC_72_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_21, data_out=>output_MAC_72_21);

	MAC_72_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_22, data_out=>output_MAC_72_22);

	MAC_72_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_23, data_out=>output_MAC_72_23);

	MAC_72_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_24, data_out=>output_MAC_72_24);

	MAC_72_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_25, data_out=>output_MAC_72_25);

	MAC_72_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_26, data_out=>output_MAC_72_26);

	MAC_72_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_27, data_out=>output_MAC_72_27);

	MAC_72_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_28, data_out=>output_MAC_72_28);

	MAC_72_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_29, data_out=>output_MAC_72_29);

	MAC_72_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_30, data_out=>output_MAC_72_30);

	MAC_72_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_72, data_in_B=>reg_input_col_31, data_out=>output_MAC_72_31);

	MAC_73_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_0, data_out=>output_MAC_73_0);

	MAC_73_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_1, data_out=>output_MAC_73_1);

	MAC_73_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_2, data_out=>output_MAC_73_2);

	MAC_73_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_3, data_out=>output_MAC_73_3);

	MAC_73_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_4, data_out=>output_MAC_73_4);

	MAC_73_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_5, data_out=>output_MAC_73_5);

	MAC_73_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_6, data_out=>output_MAC_73_6);

	MAC_73_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_7, data_out=>output_MAC_73_7);

	MAC_73_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_8, data_out=>output_MAC_73_8);

	MAC_73_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_9, data_out=>output_MAC_73_9);

	MAC_73_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_10, data_out=>output_MAC_73_10);

	MAC_73_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_11, data_out=>output_MAC_73_11);

	MAC_73_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_12, data_out=>output_MAC_73_12);

	MAC_73_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_13, data_out=>output_MAC_73_13);

	MAC_73_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_14, data_out=>output_MAC_73_14);

	MAC_73_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_15, data_out=>output_MAC_73_15);

	MAC_73_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_16, data_out=>output_MAC_73_16);

	MAC_73_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_17, data_out=>output_MAC_73_17);

	MAC_73_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_18, data_out=>output_MAC_73_18);

	MAC_73_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_19, data_out=>output_MAC_73_19);

	MAC_73_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_20, data_out=>output_MAC_73_20);

	MAC_73_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_21, data_out=>output_MAC_73_21);

	MAC_73_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_22, data_out=>output_MAC_73_22);

	MAC_73_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_23, data_out=>output_MAC_73_23);

	MAC_73_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_24, data_out=>output_MAC_73_24);

	MAC_73_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_25, data_out=>output_MAC_73_25);

	MAC_73_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_26, data_out=>output_MAC_73_26);

	MAC_73_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_27, data_out=>output_MAC_73_27);

	MAC_73_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_28, data_out=>output_MAC_73_28);

	MAC_73_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_29, data_out=>output_MAC_73_29);

	MAC_73_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_30, data_out=>output_MAC_73_30);

	MAC_73_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_73, data_in_B=>reg_input_col_31, data_out=>output_MAC_73_31);

	MAC_74_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_0, data_out=>output_MAC_74_0);

	MAC_74_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_1, data_out=>output_MAC_74_1);

	MAC_74_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_2, data_out=>output_MAC_74_2);

	MAC_74_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_3, data_out=>output_MAC_74_3);

	MAC_74_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_4, data_out=>output_MAC_74_4);

	MAC_74_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_5, data_out=>output_MAC_74_5);

	MAC_74_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_6, data_out=>output_MAC_74_6);

	MAC_74_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_7, data_out=>output_MAC_74_7);

	MAC_74_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_8, data_out=>output_MAC_74_8);

	MAC_74_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_9, data_out=>output_MAC_74_9);

	MAC_74_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_10, data_out=>output_MAC_74_10);

	MAC_74_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_11, data_out=>output_MAC_74_11);

	MAC_74_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_12, data_out=>output_MAC_74_12);

	MAC_74_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_13, data_out=>output_MAC_74_13);

	MAC_74_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_14, data_out=>output_MAC_74_14);

	MAC_74_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_15, data_out=>output_MAC_74_15);

	MAC_74_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_16, data_out=>output_MAC_74_16);

	MAC_74_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_17, data_out=>output_MAC_74_17);

	MAC_74_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_18, data_out=>output_MAC_74_18);

	MAC_74_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_19, data_out=>output_MAC_74_19);

	MAC_74_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_20, data_out=>output_MAC_74_20);

	MAC_74_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_21, data_out=>output_MAC_74_21);

	MAC_74_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_22, data_out=>output_MAC_74_22);

	MAC_74_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_23, data_out=>output_MAC_74_23);

	MAC_74_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_24, data_out=>output_MAC_74_24);

	MAC_74_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_25, data_out=>output_MAC_74_25);

	MAC_74_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_26, data_out=>output_MAC_74_26);

	MAC_74_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_27, data_out=>output_MAC_74_27);

	MAC_74_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_28, data_out=>output_MAC_74_28);

	MAC_74_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_29, data_out=>output_MAC_74_29);

	MAC_74_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_30, data_out=>output_MAC_74_30);

	MAC_74_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_74, data_in_B=>reg_input_col_31, data_out=>output_MAC_74_31);

	MAC_75_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_0, data_out=>output_MAC_75_0);

	MAC_75_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_1, data_out=>output_MAC_75_1);

	MAC_75_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_2, data_out=>output_MAC_75_2);

	MAC_75_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_3, data_out=>output_MAC_75_3);

	MAC_75_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_4, data_out=>output_MAC_75_4);

	MAC_75_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_5, data_out=>output_MAC_75_5);

	MAC_75_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_6, data_out=>output_MAC_75_6);

	MAC_75_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_7, data_out=>output_MAC_75_7);

	MAC_75_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_8, data_out=>output_MAC_75_8);

	MAC_75_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_9, data_out=>output_MAC_75_9);

	MAC_75_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_10, data_out=>output_MAC_75_10);

	MAC_75_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_11, data_out=>output_MAC_75_11);

	MAC_75_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_12, data_out=>output_MAC_75_12);

	MAC_75_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_13, data_out=>output_MAC_75_13);

	MAC_75_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_14, data_out=>output_MAC_75_14);

	MAC_75_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_15, data_out=>output_MAC_75_15);

	MAC_75_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_16, data_out=>output_MAC_75_16);

	MAC_75_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_17, data_out=>output_MAC_75_17);

	MAC_75_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_18, data_out=>output_MAC_75_18);

	MAC_75_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_19, data_out=>output_MAC_75_19);

	MAC_75_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_20, data_out=>output_MAC_75_20);

	MAC_75_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_21, data_out=>output_MAC_75_21);

	MAC_75_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_22, data_out=>output_MAC_75_22);

	MAC_75_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_23, data_out=>output_MAC_75_23);

	MAC_75_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_24, data_out=>output_MAC_75_24);

	MAC_75_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_25, data_out=>output_MAC_75_25);

	MAC_75_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_26, data_out=>output_MAC_75_26);

	MAC_75_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_27, data_out=>output_MAC_75_27);

	MAC_75_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_28, data_out=>output_MAC_75_28);

	MAC_75_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_29, data_out=>output_MAC_75_29);

	MAC_75_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_30, data_out=>output_MAC_75_30);

	MAC_75_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_75, data_in_B=>reg_input_col_31, data_out=>output_MAC_75_31);

	MAC_76_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_0, data_out=>output_MAC_76_0);

	MAC_76_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_1, data_out=>output_MAC_76_1);

	MAC_76_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_2, data_out=>output_MAC_76_2);

	MAC_76_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_3, data_out=>output_MAC_76_3);

	MAC_76_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_4, data_out=>output_MAC_76_4);

	MAC_76_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_5, data_out=>output_MAC_76_5);

	MAC_76_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_6, data_out=>output_MAC_76_6);

	MAC_76_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_7, data_out=>output_MAC_76_7);

	MAC_76_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_8, data_out=>output_MAC_76_8);

	MAC_76_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_9, data_out=>output_MAC_76_9);

	MAC_76_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_10, data_out=>output_MAC_76_10);

	MAC_76_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_11, data_out=>output_MAC_76_11);

	MAC_76_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_12, data_out=>output_MAC_76_12);

	MAC_76_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_13, data_out=>output_MAC_76_13);

	MAC_76_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_14, data_out=>output_MAC_76_14);

	MAC_76_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_15, data_out=>output_MAC_76_15);

	MAC_76_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_16, data_out=>output_MAC_76_16);

	MAC_76_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_17, data_out=>output_MAC_76_17);

	MAC_76_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_18, data_out=>output_MAC_76_18);

	MAC_76_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_19, data_out=>output_MAC_76_19);

	MAC_76_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_20, data_out=>output_MAC_76_20);

	MAC_76_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_21, data_out=>output_MAC_76_21);

	MAC_76_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_22, data_out=>output_MAC_76_22);

	MAC_76_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_23, data_out=>output_MAC_76_23);

	MAC_76_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_24, data_out=>output_MAC_76_24);

	MAC_76_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_25, data_out=>output_MAC_76_25);

	MAC_76_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_26, data_out=>output_MAC_76_26);

	MAC_76_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_27, data_out=>output_MAC_76_27);

	MAC_76_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_28, data_out=>output_MAC_76_28);

	MAC_76_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_29, data_out=>output_MAC_76_29);

	MAC_76_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_30, data_out=>output_MAC_76_30);

	MAC_76_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_76, data_in_B=>reg_input_col_31, data_out=>output_MAC_76_31);

	MAC_77_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_0, data_out=>output_MAC_77_0);

	MAC_77_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_1, data_out=>output_MAC_77_1);

	MAC_77_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_2, data_out=>output_MAC_77_2);

	MAC_77_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_3, data_out=>output_MAC_77_3);

	MAC_77_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_4, data_out=>output_MAC_77_4);

	MAC_77_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_5, data_out=>output_MAC_77_5);

	MAC_77_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_6, data_out=>output_MAC_77_6);

	MAC_77_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_7, data_out=>output_MAC_77_7);

	MAC_77_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_8, data_out=>output_MAC_77_8);

	MAC_77_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_9, data_out=>output_MAC_77_9);

	MAC_77_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_10, data_out=>output_MAC_77_10);

	MAC_77_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_11, data_out=>output_MAC_77_11);

	MAC_77_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_12, data_out=>output_MAC_77_12);

	MAC_77_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_13, data_out=>output_MAC_77_13);

	MAC_77_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_14, data_out=>output_MAC_77_14);

	MAC_77_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_15, data_out=>output_MAC_77_15);

	MAC_77_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_16, data_out=>output_MAC_77_16);

	MAC_77_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_17, data_out=>output_MAC_77_17);

	MAC_77_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_18, data_out=>output_MAC_77_18);

	MAC_77_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_19, data_out=>output_MAC_77_19);

	MAC_77_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_20, data_out=>output_MAC_77_20);

	MAC_77_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_21, data_out=>output_MAC_77_21);

	MAC_77_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_22, data_out=>output_MAC_77_22);

	MAC_77_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_23, data_out=>output_MAC_77_23);

	MAC_77_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_24, data_out=>output_MAC_77_24);

	MAC_77_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_25, data_out=>output_MAC_77_25);

	MAC_77_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_26, data_out=>output_MAC_77_26);

	MAC_77_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_27, data_out=>output_MAC_77_27);

	MAC_77_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_28, data_out=>output_MAC_77_28);

	MAC_77_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_29, data_out=>output_MAC_77_29);

	MAC_77_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_30, data_out=>output_MAC_77_30);

	MAC_77_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_77, data_in_B=>reg_input_col_31, data_out=>output_MAC_77_31);

	MAC_78_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_0, data_out=>output_MAC_78_0);

	MAC_78_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_1, data_out=>output_MAC_78_1);

	MAC_78_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_2, data_out=>output_MAC_78_2);

	MAC_78_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_3, data_out=>output_MAC_78_3);

	MAC_78_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_4, data_out=>output_MAC_78_4);

	MAC_78_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_5, data_out=>output_MAC_78_5);

	MAC_78_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_6, data_out=>output_MAC_78_6);

	MAC_78_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_7, data_out=>output_MAC_78_7);

	MAC_78_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_8, data_out=>output_MAC_78_8);

	MAC_78_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_9, data_out=>output_MAC_78_9);

	MAC_78_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_10, data_out=>output_MAC_78_10);

	MAC_78_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_11, data_out=>output_MAC_78_11);

	MAC_78_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_12, data_out=>output_MAC_78_12);

	MAC_78_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_13, data_out=>output_MAC_78_13);

	MAC_78_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_14, data_out=>output_MAC_78_14);

	MAC_78_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_15, data_out=>output_MAC_78_15);

	MAC_78_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_16, data_out=>output_MAC_78_16);

	MAC_78_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_17, data_out=>output_MAC_78_17);

	MAC_78_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_18, data_out=>output_MAC_78_18);

	MAC_78_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_19, data_out=>output_MAC_78_19);

	MAC_78_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_20, data_out=>output_MAC_78_20);

	MAC_78_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_21, data_out=>output_MAC_78_21);

	MAC_78_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_22, data_out=>output_MAC_78_22);

	MAC_78_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_23, data_out=>output_MAC_78_23);

	MAC_78_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_24, data_out=>output_MAC_78_24);

	MAC_78_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_25, data_out=>output_MAC_78_25);

	MAC_78_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_26, data_out=>output_MAC_78_26);

	MAC_78_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_27, data_out=>output_MAC_78_27);

	MAC_78_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_28, data_out=>output_MAC_78_28);

	MAC_78_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_29, data_out=>output_MAC_78_29);

	MAC_78_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_30, data_out=>output_MAC_78_30);

	MAC_78_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_78, data_in_B=>reg_input_col_31, data_out=>output_MAC_78_31);

	MAC_79_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_0, data_out=>output_MAC_79_0);

	MAC_79_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_1, data_out=>output_MAC_79_1);

	MAC_79_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_2, data_out=>output_MAC_79_2);

	MAC_79_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_3, data_out=>output_MAC_79_3);

	MAC_79_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_4, data_out=>output_MAC_79_4);

	MAC_79_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_5, data_out=>output_MAC_79_5);

	MAC_79_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_6, data_out=>output_MAC_79_6);

	MAC_79_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_7, data_out=>output_MAC_79_7);

	MAC_79_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_8, data_out=>output_MAC_79_8);

	MAC_79_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_9, data_out=>output_MAC_79_9);

	MAC_79_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_10, data_out=>output_MAC_79_10);

	MAC_79_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_11, data_out=>output_MAC_79_11);

	MAC_79_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_12, data_out=>output_MAC_79_12);

	MAC_79_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_13, data_out=>output_MAC_79_13);

	MAC_79_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_14, data_out=>output_MAC_79_14);

	MAC_79_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_15, data_out=>output_MAC_79_15);

	MAC_79_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_16, data_out=>output_MAC_79_16);

	MAC_79_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_17, data_out=>output_MAC_79_17);

	MAC_79_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_18, data_out=>output_MAC_79_18);

	MAC_79_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_19, data_out=>output_MAC_79_19);

	MAC_79_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_20, data_out=>output_MAC_79_20);

	MAC_79_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_21, data_out=>output_MAC_79_21);

	MAC_79_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_22, data_out=>output_MAC_79_22);

	MAC_79_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_23, data_out=>output_MAC_79_23);

	MAC_79_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_24, data_out=>output_MAC_79_24);

	MAC_79_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_25, data_out=>output_MAC_79_25);

	MAC_79_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_26, data_out=>output_MAC_79_26);

	MAC_79_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_27, data_out=>output_MAC_79_27);

	MAC_79_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_28, data_out=>output_MAC_79_28);

	MAC_79_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_29, data_out=>output_MAC_79_29);

	MAC_79_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_30, data_out=>output_MAC_79_30);

	MAC_79_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_79, data_in_B=>reg_input_col_31, data_out=>output_MAC_79_31);

	MAC_80_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_0, data_out=>output_MAC_80_0);

	MAC_80_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_1, data_out=>output_MAC_80_1);

	MAC_80_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_2, data_out=>output_MAC_80_2);

	MAC_80_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_3, data_out=>output_MAC_80_3);

	MAC_80_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_4, data_out=>output_MAC_80_4);

	MAC_80_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_5, data_out=>output_MAC_80_5);

	MAC_80_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_6, data_out=>output_MAC_80_6);

	MAC_80_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_7, data_out=>output_MAC_80_7);

	MAC_80_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_8, data_out=>output_MAC_80_8);

	MAC_80_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_9, data_out=>output_MAC_80_9);

	MAC_80_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_10, data_out=>output_MAC_80_10);

	MAC_80_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_11, data_out=>output_MAC_80_11);

	MAC_80_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_12, data_out=>output_MAC_80_12);

	MAC_80_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_13, data_out=>output_MAC_80_13);

	MAC_80_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_14, data_out=>output_MAC_80_14);

	MAC_80_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_15, data_out=>output_MAC_80_15);

	MAC_80_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_16, data_out=>output_MAC_80_16);

	MAC_80_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_17, data_out=>output_MAC_80_17);

	MAC_80_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_18, data_out=>output_MAC_80_18);

	MAC_80_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_19, data_out=>output_MAC_80_19);

	MAC_80_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_20, data_out=>output_MAC_80_20);

	MAC_80_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_21, data_out=>output_MAC_80_21);

	MAC_80_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_22, data_out=>output_MAC_80_22);

	MAC_80_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_23, data_out=>output_MAC_80_23);

	MAC_80_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_24, data_out=>output_MAC_80_24);

	MAC_80_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_25, data_out=>output_MAC_80_25);

	MAC_80_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_26, data_out=>output_MAC_80_26);

	MAC_80_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_27, data_out=>output_MAC_80_27);

	MAC_80_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_28, data_out=>output_MAC_80_28);

	MAC_80_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_29, data_out=>output_MAC_80_29);

	MAC_80_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_30, data_out=>output_MAC_80_30);

	MAC_80_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_80, data_in_B=>reg_input_col_31, data_out=>output_MAC_80_31);

	MAC_81_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_0, data_out=>output_MAC_81_0);

	MAC_81_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_1, data_out=>output_MAC_81_1);

	MAC_81_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_2, data_out=>output_MAC_81_2);

	MAC_81_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_3, data_out=>output_MAC_81_3);

	MAC_81_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_4, data_out=>output_MAC_81_4);

	MAC_81_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_5, data_out=>output_MAC_81_5);

	MAC_81_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_6, data_out=>output_MAC_81_6);

	MAC_81_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_7, data_out=>output_MAC_81_7);

	MAC_81_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_8, data_out=>output_MAC_81_8);

	MAC_81_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_9, data_out=>output_MAC_81_9);

	MAC_81_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_10, data_out=>output_MAC_81_10);

	MAC_81_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_11, data_out=>output_MAC_81_11);

	MAC_81_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_12, data_out=>output_MAC_81_12);

	MAC_81_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_13, data_out=>output_MAC_81_13);

	MAC_81_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_14, data_out=>output_MAC_81_14);

	MAC_81_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_15, data_out=>output_MAC_81_15);

	MAC_81_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_16, data_out=>output_MAC_81_16);

	MAC_81_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_17, data_out=>output_MAC_81_17);

	MAC_81_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_18, data_out=>output_MAC_81_18);

	MAC_81_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_19, data_out=>output_MAC_81_19);

	MAC_81_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_20, data_out=>output_MAC_81_20);

	MAC_81_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_21, data_out=>output_MAC_81_21);

	MAC_81_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_22, data_out=>output_MAC_81_22);

	MAC_81_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_23, data_out=>output_MAC_81_23);

	MAC_81_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_24, data_out=>output_MAC_81_24);

	MAC_81_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_25, data_out=>output_MAC_81_25);

	MAC_81_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_26, data_out=>output_MAC_81_26);

	MAC_81_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_27, data_out=>output_MAC_81_27);

	MAC_81_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_28, data_out=>output_MAC_81_28);

	MAC_81_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_29, data_out=>output_MAC_81_29);

	MAC_81_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_30, data_out=>output_MAC_81_30);

	MAC_81_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_81, data_in_B=>reg_input_col_31, data_out=>output_MAC_81_31);

	MAC_82_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_0, data_out=>output_MAC_82_0);

	MAC_82_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_1, data_out=>output_MAC_82_1);

	MAC_82_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_2, data_out=>output_MAC_82_2);

	MAC_82_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_3, data_out=>output_MAC_82_3);

	MAC_82_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_4, data_out=>output_MAC_82_4);

	MAC_82_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_5, data_out=>output_MAC_82_5);

	MAC_82_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_6, data_out=>output_MAC_82_6);

	MAC_82_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_7, data_out=>output_MAC_82_7);

	MAC_82_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_8, data_out=>output_MAC_82_8);

	MAC_82_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_9, data_out=>output_MAC_82_9);

	MAC_82_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_10, data_out=>output_MAC_82_10);

	MAC_82_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_11, data_out=>output_MAC_82_11);

	MAC_82_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_12, data_out=>output_MAC_82_12);

	MAC_82_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_13, data_out=>output_MAC_82_13);

	MAC_82_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_14, data_out=>output_MAC_82_14);

	MAC_82_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_15, data_out=>output_MAC_82_15);

	MAC_82_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_16, data_out=>output_MAC_82_16);

	MAC_82_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_17, data_out=>output_MAC_82_17);

	MAC_82_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_18, data_out=>output_MAC_82_18);

	MAC_82_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_19, data_out=>output_MAC_82_19);

	MAC_82_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_20, data_out=>output_MAC_82_20);

	MAC_82_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_21, data_out=>output_MAC_82_21);

	MAC_82_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_22, data_out=>output_MAC_82_22);

	MAC_82_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_23, data_out=>output_MAC_82_23);

	MAC_82_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_24, data_out=>output_MAC_82_24);

	MAC_82_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_25, data_out=>output_MAC_82_25);

	MAC_82_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_26, data_out=>output_MAC_82_26);

	MAC_82_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_27, data_out=>output_MAC_82_27);

	MAC_82_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_28, data_out=>output_MAC_82_28);

	MAC_82_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_29, data_out=>output_MAC_82_29);

	MAC_82_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_30, data_out=>output_MAC_82_30);

	MAC_82_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_82, data_in_B=>reg_input_col_31, data_out=>output_MAC_82_31);

	MAC_83_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_0, data_out=>output_MAC_83_0);

	MAC_83_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_1, data_out=>output_MAC_83_1);

	MAC_83_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_2, data_out=>output_MAC_83_2);

	MAC_83_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_3, data_out=>output_MAC_83_3);

	MAC_83_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_4, data_out=>output_MAC_83_4);

	MAC_83_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_5, data_out=>output_MAC_83_5);

	MAC_83_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_6, data_out=>output_MAC_83_6);

	MAC_83_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_7, data_out=>output_MAC_83_7);

	MAC_83_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_8, data_out=>output_MAC_83_8);

	MAC_83_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_9, data_out=>output_MAC_83_9);

	MAC_83_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_10, data_out=>output_MAC_83_10);

	MAC_83_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_11, data_out=>output_MAC_83_11);

	MAC_83_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_12, data_out=>output_MAC_83_12);

	MAC_83_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_13, data_out=>output_MAC_83_13);

	MAC_83_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_14, data_out=>output_MAC_83_14);

	MAC_83_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_15, data_out=>output_MAC_83_15);

	MAC_83_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_16, data_out=>output_MAC_83_16);

	MAC_83_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_17, data_out=>output_MAC_83_17);

	MAC_83_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_18, data_out=>output_MAC_83_18);

	MAC_83_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_19, data_out=>output_MAC_83_19);

	MAC_83_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_20, data_out=>output_MAC_83_20);

	MAC_83_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_21, data_out=>output_MAC_83_21);

	MAC_83_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_22, data_out=>output_MAC_83_22);

	MAC_83_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_23, data_out=>output_MAC_83_23);

	MAC_83_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_24, data_out=>output_MAC_83_24);

	MAC_83_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_25, data_out=>output_MAC_83_25);

	MAC_83_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_26, data_out=>output_MAC_83_26);

	MAC_83_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_27, data_out=>output_MAC_83_27);

	MAC_83_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_28, data_out=>output_MAC_83_28);

	MAC_83_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_29, data_out=>output_MAC_83_29);

	MAC_83_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_30, data_out=>output_MAC_83_30);

	MAC_83_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_83, data_in_B=>reg_input_col_31, data_out=>output_MAC_83_31);

	MAC_84_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_0, data_out=>output_MAC_84_0);

	MAC_84_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_1, data_out=>output_MAC_84_1);

	MAC_84_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_2, data_out=>output_MAC_84_2);

	MAC_84_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_3, data_out=>output_MAC_84_3);

	MAC_84_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_4, data_out=>output_MAC_84_4);

	MAC_84_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_5, data_out=>output_MAC_84_5);

	MAC_84_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_6, data_out=>output_MAC_84_6);

	MAC_84_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_7, data_out=>output_MAC_84_7);

	MAC_84_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_8, data_out=>output_MAC_84_8);

	MAC_84_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_9, data_out=>output_MAC_84_9);

	MAC_84_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_10, data_out=>output_MAC_84_10);

	MAC_84_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_11, data_out=>output_MAC_84_11);

	MAC_84_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_12, data_out=>output_MAC_84_12);

	MAC_84_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_13, data_out=>output_MAC_84_13);

	MAC_84_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_14, data_out=>output_MAC_84_14);

	MAC_84_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_15, data_out=>output_MAC_84_15);

	MAC_84_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_16, data_out=>output_MAC_84_16);

	MAC_84_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_17, data_out=>output_MAC_84_17);

	MAC_84_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_18, data_out=>output_MAC_84_18);

	MAC_84_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_19, data_out=>output_MAC_84_19);

	MAC_84_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_20, data_out=>output_MAC_84_20);

	MAC_84_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_21, data_out=>output_MAC_84_21);

	MAC_84_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_22, data_out=>output_MAC_84_22);

	MAC_84_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_23, data_out=>output_MAC_84_23);

	MAC_84_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_24, data_out=>output_MAC_84_24);

	MAC_84_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_25, data_out=>output_MAC_84_25);

	MAC_84_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_26, data_out=>output_MAC_84_26);

	MAC_84_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_27, data_out=>output_MAC_84_27);

	MAC_84_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_28, data_out=>output_MAC_84_28);

	MAC_84_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_29, data_out=>output_MAC_84_29);

	MAC_84_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_30, data_out=>output_MAC_84_30);

	MAC_84_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_84, data_in_B=>reg_input_col_31, data_out=>output_MAC_84_31);

	MAC_85_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_0, data_out=>output_MAC_85_0);

	MAC_85_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_1, data_out=>output_MAC_85_1);

	MAC_85_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_2, data_out=>output_MAC_85_2);

	MAC_85_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_3, data_out=>output_MAC_85_3);

	MAC_85_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_4, data_out=>output_MAC_85_4);

	MAC_85_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_5, data_out=>output_MAC_85_5);

	MAC_85_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_6, data_out=>output_MAC_85_6);

	MAC_85_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_7, data_out=>output_MAC_85_7);

	MAC_85_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_8, data_out=>output_MAC_85_8);

	MAC_85_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_9, data_out=>output_MAC_85_9);

	MAC_85_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_10, data_out=>output_MAC_85_10);

	MAC_85_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_11, data_out=>output_MAC_85_11);

	MAC_85_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_12, data_out=>output_MAC_85_12);

	MAC_85_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_13, data_out=>output_MAC_85_13);

	MAC_85_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_14, data_out=>output_MAC_85_14);

	MAC_85_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_15, data_out=>output_MAC_85_15);

	MAC_85_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_16, data_out=>output_MAC_85_16);

	MAC_85_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_17, data_out=>output_MAC_85_17);

	MAC_85_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_18, data_out=>output_MAC_85_18);

	MAC_85_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_19, data_out=>output_MAC_85_19);

	MAC_85_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_20, data_out=>output_MAC_85_20);

	MAC_85_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_21, data_out=>output_MAC_85_21);

	MAC_85_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_22, data_out=>output_MAC_85_22);

	MAC_85_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_23, data_out=>output_MAC_85_23);

	MAC_85_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_24, data_out=>output_MAC_85_24);

	MAC_85_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_25, data_out=>output_MAC_85_25);

	MAC_85_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_26, data_out=>output_MAC_85_26);

	MAC_85_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_27, data_out=>output_MAC_85_27);

	MAC_85_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_28, data_out=>output_MAC_85_28);

	MAC_85_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_29, data_out=>output_MAC_85_29);

	MAC_85_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_30, data_out=>output_MAC_85_30);

	MAC_85_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_85, data_in_B=>reg_input_col_31, data_out=>output_MAC_85_31);

	MAC_86_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_0, data_out=>output_MAC_86_0);

	MAC_86_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_1, data_out=>output_MAC_86_1);

	MAC_86_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_2, data_out=>output_MAC_86_2);

	MAC_86_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_3, data_out=>output_MAC_86_3);

	MAC_86_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_4, data_out=>output_MAC_86_4);

	MAC_86_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_5, data_out=>output_MAC_86_5);

	MAC_86_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_6, data_out=>output_MAC_86_6);

	MAC_86_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_7, data_out=>output_MAC_86_7);

	MAC_86_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_8, data_out=>output_MAC_86_8);

	MAC_86_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_9, data_out=>output_MAC_86_9);

	MAC_86_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_10, data_out=>output_MAC_86_10);

	MAC_86_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_11, data_out=>output_MAC_86_11);

	MAC_86_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_12, data_out=>output_MAC_86_12);

	MAC_86_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_13, data_out=>output_MAC_86_13);

	MAC_86_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_14, data_out=>output_MAC_86_14);

	MAC_86_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_15, data_out=>output_MAC_86_15);

	MAC_86_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_16, data_out=>output_MAC_86_16);

	MAC_86_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_17, data_out=>output_MAC_86_17);

	MAC_86_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_18, data_out=>output_MAC_86_18);

	MAC_86_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_19, data_out=>output_MAC_86_19);

	MAC_86_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_20, data_out=>output_MAC_86_20);

	MAC_86_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_21, data_out=>output_MAC_86_21);

	MAC_86_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_22, data_out=>output_MAC_86_22);

	MAC_86_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_23, data_out=>output_MAC_86_23);

	MAC_86_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_24, data_out=>output_MAC_86_24);

	MAC_86_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_25, data_out=>output_MAC_86_25);

	MAC_86_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_26, data_out=>output_MAC_86_26);

	MAC_86_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_27, data_out=>output_MAC_86_27);

	MAC_86_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_28, data_out=>output_MAC_86_28);

	MAC_86_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_29, data_out=>output_MAC_86_29);

	MAC_86_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_30, data_out=>output_MAC_86_30);

	MAC_86_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_86, data_in_B=>reg_input_col_31, data_out=>output_MAC_86_31);

	MAC_87_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_0, data_out=>output_MAC_87_0);

	MAC_87_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_1, data_out=>output_MAC_87_1);

	MAC_87_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_2, data_out=>output_MAC_87_2);

	MAC_87_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_3, data_out=>output_MAC_87_3);

	MAC_87_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_4, data_out=>output_MAC_87_4);

	MAC_87_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_5, data_out=>output_MAC_87_5);

	MAC_87_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_6, data_out=>output_MAC_87_6);

	MAC_87_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_7, data_out=>output_MAC_87_7);

	MAC_87_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_8, data_out=>output_MAC_87_8);

	MAC_87_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_9, data_out=>output_MAC_87_9);

	MAC_87_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_10, data_out=>output_MAC_87_10);

	MAC_87_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_11, data_out=>output_MAC_87_11);

	MAC_87_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_12, data_out=>output_MAC_87_12);

	MAC_87_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_13, data_out=>output_MAC_87_13);

	MAC_87_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_14, data_out=>output_MAC_87_14);

	MAC_87_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_15, data_out=>output_MAC_87_15);

	MAC_87_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_16, data_out=>output_MAC_87_16);

	MAC_87_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_17, data_out=>output_MAC_87_17);

	MAC_87_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_18, data_out=>output_MAC_87_18);

	MAC_87_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_19, data_out=>output_MAC_87_19);

	MAC_87_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_20, data_out=>output_MAC_87_20);

	MAC_87_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_21, data_out=>output_MAC_87_21);

	MAC_87_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_22, data_out=>output_MAC_87_22);

	MAC_87_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_23, data_out=>output_MAC_87_23);

	MAC_87_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_24, data_out=>output_MAC_87_24);

	MAC_87_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_25, data_out=>output_MAC_87_25);

	MAC_87_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_26, data_out=>output_MAC_87_26);

	MAC_87_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_27, data_out=>output_MAC_87_27);

	MAC_87_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_28, data_out=>output_MAC_87_28);

	MAC_87_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_29, data_out=>output_MAC_87_29);

	MAC_87_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_30, data_out=>output_MAC_87_30);

	MAC_87_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_87, data_in_B=>reg_input_col_31, data_out=>output_MAC_87_31);

	MAC_88_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_0, data_out=>output_MAC_88_0);

	MAC_88_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_1, data_out=>output_MAC_88_1);

	MAC_88_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_2, data_out=>output_MAC_88_2);

	MAC_88_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_3, data_out=>output_MAC_88_3);

	MAC_88_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_4, data_out=>output_MAC_88_4);

	MAC_88_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_5, data_out=>output_MAC_88_5);

	MAC_88_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_6, data_out=>output_MAC_88_6);

	MAC_88_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_7, data_out=>output_MAC_88_7);

	MAC_88_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_8, data_out=>output_MAC_88_8);

	MAC_88_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_9, data_out=>output_MAC_88_9);

	MAC_88_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_10, data_out=>output_MAC_88_10);

	MAC_88_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_11, data_out=>output_MAC_88_11);

	MAC_88_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_12, data_out=>output_MAC_88_12);

	MAC_88_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_13, data_out=>output_MAC_88_13);

	MAC_88_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_14, data_out=>output_MAC_88_14);

	MAC_88_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_15, data_out=>output_MAC_88_15);

	MAC_88_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_16, data_out=>output_MAC_88_16);

	MAC_88_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_17, data_out=>output_MAC_88_17);

	MAC_88_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_18, data_out=>output_MAC_88_18);

	MAC_88_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_19, data_out=>output_MAC_88_19);

	MAC_88_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_20, data_out=>output_MAC_88_20);

	MAC_88_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_21, data_out=>output_MAC_88_21);

	MAC_88_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_22, data_out=>output_MAC_88_22);

	MAC_88_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_23, data_out=>output_MAC_88_23);

	MAC_88_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_24, data_out=>output_MAC_88_24);

	MAC_88_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_25, data_out=>output_MAC_88_25);

	MAC_88_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_26, data_out=>output_MAC_88_26);

	MAC_88_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_27, data_out=>output_MAC_88_27);

	MAC_88_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_28, data_out=>output_MAC_88_28);

	MAC_88_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_29, data_out=>output_MAC_88_29);

	MAC_88_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_30, data_out=>output_MAC_88_30);

	MAC_88_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_88, data_in_B=>reg_input_col_31, data_out=>output_MAC_88_31);

	MAC_89_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_0, data_out=>output_MAC_89_0);

	MAC_89_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_1, data_out=>output_MAC_89_1);

	MAC_89_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_2, data_out=>output_MAC_89_2);

	MAC_89_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_3, data_out=>output_MAC_89_3);

	MAC_89_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_4, data_out=>output_MAC_89_4);

	MAC_89_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_5, data_out=>output_MAC_89_5);

	MAC_89_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_6, data_out=>output_MAC_89_6);

	MAC_89_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_7, data_out=>output_MAC_89_7);

	MAC_89_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_8, data_out=>output_MAC_89_8);

	MAC_89_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_9, data_out=>output_MAC_89_9);

	MAC_89_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_10, data_out=>output_MAC_89_10);

	MAC_89_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_11, data_out=>output_MAC_89_11);

	MAC_89_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_12, data_out=>output_MAC_89_12);

	MAC_89_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_13, data_out=>output_MAC_89_13);

	MAC_89_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_14, data_out=>output_MAC_89_14);

	MAC_89_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_15, data_out=>output_MAC_89_15);

	MAC_89_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_16, data_out=>output_MAC_89_16);

	MAC_89_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_17, data_out=>output_MAC_89_17);

	MAC_89_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_18, data_out=>output_MAC_89_18);

	MAC_89_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_19, data_out=>output_MAC_89_19);

	MAC_89_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_20, data_out=>output_MAC_89_20);

	MAC_89_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_21, data_out=>output_MAC_89_21);

	MAC_89_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_22, data_out=>output_MAC_89_22);

	MAC_89_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_23, data_out=>output_MAC_89_23);

	MAC_89_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_24, data_out=>output_MAC_89_24);

	MAC_89_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_25, data_out=>output_MAC_89_25);

	MAC_89_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_26, data_out=>output_MAC_89_26);

	MAC_89_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_27, data_out=>output_MAC_89_27);

	MAC_89_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_28, data_out=>output_MAC_89_28);

	MAC_89_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_29, data_out=>output_MAC_89_29);

	MAC_89_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_30, data_out=>output_MAC_89_30);

	MAC_89_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_89, data_in_B=>reg_input_col_31, data_out=>output_MAC_89_31);

	MAC_90_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_0, data_out=>output_MAC_90_0);

	MAC_90_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_1, data_out=>output_MAC_90_1);

	MAC_90_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_2, data_out=>output_MAC_90_2);

	MAC_90_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_3, data_out=>output_MAC_90_3);

	MAC_90_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_4, data_out=>output_MAC_90_4);

	MAC_90_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_5, data_out=>output_MAC_90_5);

	MAC_90_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_6, data_out=>output_MAC_90_6);

	MAC_90_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_7, data_out=>output_MAC_90_7);

	MAC_90_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_8, data_out=>output_MAC_90_8);

	MAC_90_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_9, data_out=>output_MAC_90_9);

	MAC_90_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_10, data_out=>output_MAC_90_10);

	MAC_90_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_11, data_out=>output_MAC_90_11);

	MAC_90_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_12, data_out=>output_MAC_90_12);

	MAC_90_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_13, data_out=>output_MAC_90_13);

	MAC_90_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_14, data_out=>output_MAC_90_14);

	MAC_90_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_15, data_out=>output_MAC_90_15);

	MAC_90_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_16, data_out=>output_MAC_90_16);

	MAC_90_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_17, data_out=>output_MAC_90_17);

	MAC_90_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_18, data_out=>output_MAC_90_18);

	MAC_90_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_19, data_out=>output_MAC_90_19);

	MAC_90_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_20, data_out=>output_MAC_90_20);

	MAC_90_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_21, data_out=>output_MAC_90_21);

	MAC_90_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_22, data_out=>output_MAC_90_22);

	MAC_90_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_23, data_out=>output_MAC_90_23);

	MAC_90_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_24, data_out=>output_MAC_90_24);

	MAC_90_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_25, data_out=>output_MAC_90_25);

	MAC_90_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_26, data_out=>output_MAC_90_26);

	MAC_90_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_27, data_out=>output_MAC_90_27);

	MAC_90_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_28, data_out=>output_MAC_90_28);

	MAC_90_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_29, data_out=>output_MAC_90_29);

	MAC_90_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_30, data_out=>output_MAC_90_30);

	MAC_90_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_90, data_in_B=>reg_input_col_31, data_out=>output_MAC_90_31);

	MAC_91_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_0, data_out=>output_MAC_91_0);

	MAC_91_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_1, data_out=>output_MAC_91_1);

	MAC_91_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_2, data_out=>output_MAC_91_2);

	MAC_91_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_3, data_out=>output_MAC_91_3);

	MAC_91_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_4, data_out=>output_MAC_91_4);

	MAC_91_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_5, data_out=>output_MAC_91_5);

	MAC_91_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_6, data_out=>output_MAC_91_6);

	MAC_91_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_7, data_out=>output_MAC_91_7);

	MAC_91_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_8, data_out=>output_MAC_91_8);

	MAC_91_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_9, data_out=>output_MAC_91_9);

	MAC_91_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_10, data_out=>output_MAC_91_10);

	MAC_91_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_11, data_out=>output_MAC_91_11);

	MAC_91_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_12, data_out=>output_MAC_91_12);

	MAC_91_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_13, data_out=>output_MAC_91_13);

	MAC_91_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_14, data_out=>output_MAC_91_14);

	MAC_91_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_15, data_out=>output_MAC_91_15);

	MAC_91_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_16, data_out=>output_MAC_91_16);

	MAC_91_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_17, data_out=>output_MAC_91_17);

	MAC_91_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_18, data_out=>output_MAC_91_18);

	MAC_91_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_19, data_out=>output_MAC_91_19);

	MAC_91_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_20, data_out=>output_MAC_91_20);

	MAC_91_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_21, data_out=>output_MAC_91_21);

	MAC_91_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_22, data_out=>output_MAC_91_22);

	MAC_91_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_23, data_out=>output_MAC_91_23);

	MAC_91_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_24, data_out=>output_MAC_91_24);

	MAC_91_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_25, data_out=>output_MAC_91_25);

	MAC_91_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_26, data_out=>output_MAC_91_26);

	MAC_91_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_27, data_out=>output_MAC_91_27);

	MAC_91_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_28, data_out=>output_MAC_91_28);

	MAC_91_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_29, data_out=>output_MAC_91_29);

	MAC_91_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_30, data_out=>output_MAC_91_30);

	MAC_91_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_91, data_in_B=>reg_input_col_31, data_out=>output_MAC_91_31);

	MAC_92_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_0, data_out=>output_MAC_92_0);

	MAC_92_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_1, data_out=>output_MAC_92_1);

	MAC_92_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_2, data_out=>output_MAC_92_2);

	MAC_92_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_3, data_out=>output_MAC_92_3);

	MAC_92_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_4, data_out=>output_MAC_92_4);

	MAC_92_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_5, data_out=>output_MAC_92_5);

	MAC_92_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_6, data_out=>output_MAC_92_6);

	MAC_92_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_7, data_out=>output_MAC_92_7);

	MAC_92_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_8, data_out=>output_MAC_92_8);

	MAC_92_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_9, data_out=>output_MAC_92_9);

	MAC_92_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_10, data_out=>output_MAC_92_10);

	MAC_92_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_11, data_out=>output_MAC_92_11);

	MAC_92_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_12, data_out=>output_MAC_92_12);

	MAC_92_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_13, data_out=>output_MAC_92_13);

	MAC_92_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_14, data_out=>output_MAC_92_14);

	MAC_92_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_15, data_out=>output_MAC_92_15);

	MAC_92_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_16, data_out=>output_MAC_92_16);

	MAC_92_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_17, data_out=>output_MAC_92_17);

	MAC_92_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_18, data_out=>output_MAC_92_18);

	MAC_92_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_19, data_out=>output_MAC_92_19);

	MAC_92_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_20, data_out=>output_MAC_92_20);

	MAC_92_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_21, data_out=>output_MAC_92_21);

	MAC_92_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_22, data_out=>output_MAC_92_22);

	MAC_92_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_23, data_out=>output_MAC_92_23);

	MAC_92_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_24, data_out=>output_MAC_92_24);

	MAC_92_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_25, data_out=>output_MAC_92_25);

	MAC_92_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_26, data_out=>output_MAC_92_26);

	MAC_92_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_27, data_out=>output_MAC_92_27);

	MAC_92_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_28, data_out=>output_MAC_92_28);

	MAC_92_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_29, data_out=>output_MAC_92_29);

	MAC_92_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_30, data_out=>output_MAC_92_30);

	MAC_92_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_92, data_in_B=>reg_input_col_31, data_out=>output_MAC_92_31);

	MAC_93_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_0, data_out=>output_MAC_93_0);

	MAC_93_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_1, data_out=>output_MAC_93_1);

	MAC_93_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_2, data_out=>output_MAC_93_2);

	MAC_93_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_3, data_out=>output_MAC_93_3);

	MAC_93_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_4, data_out=>output_MAC_93_4);

	MAC_93_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_5, data_out=>output_MAC_93_5);

	MAC_93_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_6, data_out=>output_MAC_93_6);

	MAC_93_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_7, data_out=>output_MAC_93_7);

	MAC_93_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_8, data_out=>output_MAC_93_8);

	MAC_93_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_9, data_out=>output_MAC_93_9);

	MAC_93_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_10, data_out=>output_MAC_93_10);

	MAC_93_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_11, data_out=>output_MAC_93_11);

	MAC_93_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_12, data_out=>output_MAC_93_12);

	MAC_93_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_13, data_out=>output_MAC_93_13);

	MAC_93_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_14, data_out=>output_MAC_93_14);

	MAC_93_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_15, data_out=>output_MAC_93_15);

	MAC_93_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_16, data_out=>output_MAC_93_16);

	MAC_93_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_17, data_out=>output_MAC_93_17);

	MAC_93_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_18, data_out=>output_MAC_93_18);

	MAC_93_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_19, data_out=>output_MAC_93_19);

	MAC_93_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_20, data_out=>output_MAC_93_20);

	MAC_93_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_21, data_out=>output_MAC_93_21);

	MAC_93_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_22, data_out=>output_MAC_93_22);

	MAC_93_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_23, data_out=>output_MAC_93_23);

	MAC_93_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_24, data_out=>output_MAC_93_24);

	MAC_93_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_25, data_out=>output_MAC_93_25);

	MAC_93_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_26, data_out=>output_MAC_93_26);

	MAC_93_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_27, data_out=>output_MAC_93_27);

	MAC_93_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_28, data_out=>output_MAC_93_28);

	MAC_93_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_29, data_out=>output_MAC_93_29);

	MAC_93_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_30, data_out=>output_MAC_93_30);

	MAC_93_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_93, data_in_B=>reg_input_col_31, data_out=>output_MAC_93_31);

	MAC_94_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_0, data_out=>output_MAC_94_0);

	MAC_94_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_1, data_out=>output_MAC_94_1);

	MAC_94_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_2, data_out=>output_MAC_94_2);

	MAC_94_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_3, data_out=>output_MAC_94_3);

	MAC_94_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_4, data_out=>output_MAC_94_4);

	MAC_94_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_5, data_out=>output_MAC_94_5);

	MAC_94_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_6, data_out=>output_MAC_94_6);

	MAC_94_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_7, data_out=>output_MAC_94_7);

	MAC_94_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_8, data_out=>output_MAC_94_8);

	MAC_94_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_9, data_out=>output_MAC_94_9);

	MAC_94_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_10, data_out=>output_MAC_94_10);

	MAC_94_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_11, data_out=>output_MAC_94_11);

	MAC_94_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_12, data_out=>output_MAC_94_12);

	MAC_94_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_13, data_out=>output_MAC_94_13);

	MAC_94_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_14, data_out=>output_MAC_94_14);

	MAC_94_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_15, data_out=>output_MAC_94_15);

	MAC_94_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_16, data_out=>output_MAC_94_16);

	MAC_94_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_17, data_out=>output_MAC_94_17);

	MAC_94_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_18, data_out=>output_MAC_94_18);

	MAC_94_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_19, data_out=>output_MAC_94_19);

	MAC_94_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_20, data_out=>output_MAC_94_20);

	MAC_94_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_21, data_out=>output_MAC_94_21);

	MAC_94_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_22, data_out=>output_MAC_94_22);

	MAC_94_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_23, data_out=>output_MAC_94_23);

	MAC_94_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_24, data_out=>output_MAC_94_24);

	MAC_94_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_25, data_out=>output_MAC_94_25);

	MAC_94_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_26, data_out=>output_MAC_94_26);

	MAC_94_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_27, data_out=>output_MAC_94_27);

	MAC_94_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_28, data_out=>output_MAC_94_28);

	MAC_94_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_29, data_out=>output_MAC_94_29);

	MAC_94_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_30, data_out=>output_MAC_94_30);

	MAC_94_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_94, data_in_B=>reg_input_col_31, data_out=>output_MAC_94_31);

	MAC_95_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_0, data_out=>output_MAC_95_0);

	MAC_95_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_1, data_out=>output_MAC_95_1);

	MAC_95_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_2, data_out=>output_MAC_95_2);

	MAC_95_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_3, data_out=>output_MAC_95_3);

	MAC_95_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_4, data_out=>output_MAC_95_4);

	MAC_95_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_5, data_out=>output_MAC_95_5);

	MAC_95_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_6, data_out=>output_MAC_95_6);

	MAC_95_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_7, data_out=>output_MAC_95_7);

	MAC_95_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_8, data_out=>output_MAC_95_8);

	MAC_95_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_9, data_out=>output_MAC_95_9);

	MAC_95_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_10, data_out=>output_MAC_95_10);

	MAC_95_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_11, data_out=>output_MAC_95_11);

	MAC_95_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_12, data_out=>output_MAC_95_12);

	MAC_95_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_13, data_out=>output_MAC_95_13);

	MAC_95_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_14, data_out=>output_MAC_95_14);

	MAC_95_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_15, data_out=>output_MAC_95_15);

	MAC_95_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_16, data_out=>output_MAC_95_16);

	MAC_95_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_17, data_out=>output_MAC_95_17);

	MAC_95_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_18, data_out=>output_MAC_95_18);

	MAC_95_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_19, data_out=>output_MAC_95_19);

	MAC_95_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_20, data_out=>output_MAC_95_20);

	MAC_95_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_21, data_out=>output_MAC_95_21);

	MAC_95_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_22, data_out=>output_MAC_95_22);

	MAC_95_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_23, data_out=>output_MAC_95_23);

	MAC_95_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_24, data_out=>output_MAC_95_24);

	MAC_95_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_25, data_out=>output_MAC_95_25);

	MAC_95_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_26, data_out=>output_MAC_95_26);

	MAC_95_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_27, data_out=>output_MAC_95_27);

	MAC_95_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_28, data_out=>output_MAC_95_28);

	MAC_95_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_29, data_out=>output_MAC_95_29);

	MAC_95_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_30, data_out=>output_MAC_95_30);

	MAC_95_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_95, data_in_B=>reg_input_col_31, data_out=>output_MAC_95_31);

	MAC_96_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_0, data_out=>output_MAC_96_0);

	MAC_96_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_1, data_out=>output_MAC_96_1);

	MAC_96_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_2, data_out=>output_MAC_96_2);

	MAC_96_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_3, data_out=>output_MAC_96_3);

	MAC_96_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_4, data_out=>output_MAC_96_4);

	MAC_96_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_5, data_out=>output_MAC_96_5);

	MAC_96_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_6, data_out=>output_MAC_96_6);

	MAC_96_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_7, data_out=>output_MAC_96_7);

	MAC_96_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_8, data_out=>output_MAC_96_8);

	MAC_96_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_9, data_out=>output_MAC_96_9);

	MAC_96_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_10, data_out=>output_MAC_96_10);

	MAC_96_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_11, data_out=>output_MAC_96_11);

	MAC_96_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_12, data_out=>output_MAC_96_12);

	MAC_96_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_13, data_out=>output_MAC_96_13);

	MAC_96_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_14, data_out=>output_MAC_96_14);

	MAC_96_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_15, data_out=>output_MAC_96_15);

	MAC_96_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_16, data_out=>output_MAC_96_16);

	MAC_96_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_17, data_out=>output_MAC_96_17);

	MAC_96_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_18, data_out=>output_MAC_96_18);

	MAC_96_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_19, data_out=>output_MAC_96_19);

	MAC_96_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_20, data_out=>output_MAC_96_20);

	MAC_96_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_21, data_out=>output_MAC_96_21);

	MAC_96_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_22, data_out=>output_MAC_96_22);

	MAC_96_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_23, data_out=>output_MAC_96_23);

	MAC_96_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_24, data_out=>output_MAC_96_24);

	MAC_96_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_25, data_out=>output_MAC_96_25);

	MAC_96_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_26, data_out=>output_MAC_96_26);

	MAC_96_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_27, data_out=>output_MAC_96_27);

	MAC_96_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_28, data_out=>output_MAC_96_28);

	MAC_96_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_29, data_out=>output_MAC_96_29);

	MAC_96_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_30, data_out=>output_MAC_96_30);

	MAC_96_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_96, data_in_B=>reg_input_col_31, data_out=>output_MAC_96_31);

	MAC_97_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_0, data_out=>output_MAC_97_0);

	MAC_97_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_1, data_out=>output_MAC_97_1);

	MAC_97_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_2, data_out=>output_MAC_97_2);

	MAC_97_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_3, data_out=>output_MAC_97_3);

	MAC_97_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_4, data_out=>output_MAC_97_4);

	MAC_97_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_5, data_out=>output_MAC_97_5);

	MAC_97_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_6, data_out=>output_MAC_97_6);

	MAC_97_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_7, data_out=>output_MAC_97_7);

	MAC_97_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_8, data_out=>output_MAC_97_8);

	MAC_97_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_9, data_out=>output_MAC_97_9);

	MAC_97_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_10, data_out=>output_MAC_97_10);

	MAC_97_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_11, data_out=>output_MAC_97_11);

	MAC_97_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_12, data_out=>output_MAC_97_12);

	MAC_97_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_13, data_out=>output_MAC_97_13);

	MAC_97_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_14, data_out=>output_MAC_97_14);

	MAC_97_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_15, data_out=>output_MAC_97_15);

	MAC_97_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_16, data_out=>output_MAC_97_16);

	MAC_97_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_17, data_out=>output_MAC_97_17);

	MAC_97_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_18, data_out=>output_MAC_97_18);

	MAC_97_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_19, data_out=>output_MAC_97_19);

	MAC_97_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_20, data_out=>output_MAC_97_20);

	MAC_97_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_21, data_out=>output_MAC_97_21);

	MAC_97_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_22, data_out=>output_MAC_97_22);

	MAC_97_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_23, data_out=>output_MAC_97_23);

	MAC_97_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_24, data_out=>output_MAC_97_24);

	MAC_97_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_25, data_out=>output_MAC_97_25);

	MAC_97_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_26, data_out=>output_MAC_97_26);

	MAC_97_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_27, data_out=>output_MAC_97_27);

	MAC_97_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_28, data_out=>output_MAC_97_28);

	MAC_97_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_29, data_out=>output_MAC_97_29);

	MAC_97_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_30, data_out=>output_MAC_97_30);

	MAC_97_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_97, data_in_B=>reg_input_col_31, data_out=>output_MAC_97_31);

	MAC_98_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_0, data_out=>output_MAC_98_0);

	MAC_98_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_1, data_out=>output_MAC_98_1);

	MAC_98_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_2, data_out=>output_MAC_98_2);

	MAC_98_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_3, data_out=>output_MAC_98_3);

	MAC_98_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_4, data_out=>output_MAC_98_4);

	MAC_98_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_5, data_out=>output_MAC_98_5);

	MAC_98_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_6, data_out=>output_MAC_98_6);

	MAC_98_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_7, data_out=>output_MAC_98_7);

	MAC_98_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_8, data_out=>output_MAC_98_8);

	MAC_98_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_9, data_out=>output_MAC_98_9);

	MAC_98_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_10, data_out=>output_MAC_98_10);

	MAC_98_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_11, data_out=>output_MAC_98_11);

	MAC_98_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_12, data_out=>output_MAC_98_12);

	MAC_98_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_13, data_out=>output_MAC_98_13);

	MAC_98_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_14, data_out=>output_MAC_98_14);

	MAC_98_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_15, data_out=>output_MAC_98_15);

	MAC_98_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_16, data_out=>output_MAC_98_16);

	MAC_98_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_17, data_out=>output_MAC_98_17);

	MAC_98_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_18, data_out=>output_MAC_98_18);

	MAC_98_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_19, data_out=>output_MAC_98_19);

	MAC_98_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_20, data_out=>output_MAC_98_20);

	MAC_98_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_21, data_out=>output_MAC_98_21);

	MAC_98_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_22, data_out=>output_MAC_98_22);

	MAC_98_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_23, data_out=>output_MAC_98_23);

	MAC_98_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_24, data_out=>output_MAC_98_24);

	MAC_98_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_25, data_out=>output_MAC_98_25);

	MAC_98_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_26, data_out=>output_MAC_98_26);

	MAC_98_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_27, data_out=>output_MAC_98_27);

	MAC_98_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_28, data_out=>output_MAC_98_28);

	MAC_98_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_29, data_out=>output_MAC_98_29);

	MAC_98_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_30, data_out=>output_MAC_98_30);

	MAC_98_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_98, data_in_B=>reg_input_col_31, data_out=>output_MAC_98_31);

	MAC_99_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_0, data_out=>output_MAC_99_0);

	MAC_99_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_1, data_out=>output_MAC_99_1);

	MAC_99_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_2, data_out=>output_MAC_99_2);

	MAC_99_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_3, data_out=>output_MAC_99_3);

	MAC_99_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_4, data_out=>output_MAC_99_4);

	MAC_99_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_5, data_out=>output_MAC_99_5);

	MAC_99_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_6, data_out=>output_MAC_99_6);

	MAC_99_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_7, data_out=>output_MAC_99_7);

	MAC_99_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_8, data_out=>output_MAC_99_8);

	MAC_99_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_9, data_out=>output_MAC_99_9);

	MAC_99_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_10, data_out=>output_MAC_99_10);

	MAC_99_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_11, data_out=>output_MAC_99_11);

	MAC_99_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_12, data_out=>output_MAC_99_12);

	MAC_99_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_13, data_out=>output_MAC_99_13);

	MAC_99_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_14, data_out=>output_MAC_99_14);

	MAC_99_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_15, data_out=>output_MAC_99_15);

	MAC_99_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_16, data_out=>output_MAC_99_16);

	MAC_99_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_17, data_out=>output_MAC_99_17);

	MAC_99_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_18, data_out=>output_MAC_99_18);

	MAC_99_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_19, data_out=>output_MAC_99_19);

	MAC_99_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_20, data_out=>output_MAC_99_20);

	MAC_99_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_21, data_out=>output_MAC_99_21);

	MAC_99_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_22, data_out=>output_MAC_99_22);

	MAC_99_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_23, data_out=>output_MAC_99_23);

	MAC_99_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_24, data_out=>output_MAC_99_24);

	MAC_99_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_25, data_out=>output_MAC_99_25);

	MAC_99_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_26, data_out=>output_MAC_99_26);

	MAC_99_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_27, data_out=>output_MAC_99_27);

	MAC_99_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_28, data_out=>output_MAC_99_28);

	MAC_99_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_29, data_out=>output_MAC_99_29);

	MAC_99_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_30, data_out=>output_MAC_99_30);

	MAC_99_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_99, data_in_B=>reg_input_col_31, data_out=>output_MAC_99_31);

	MAC_100_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_0, data_out=>output_MAC_100_0);

	MAC_100_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_1, data_out=>output_MAC_100_1);

	MAC_100_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_2, data_out=>output_MAC_100_2);

	MAC_100_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_3, data_out=>output_MAC_100_3);

	MAC_100_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_4, data_out=>output_MAC_100_4);

	MAC_100_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_5, data_out=>output_MAC_100_5);

	MAC_100_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_6, data_out=>output_MAC_100_6);

	MAC_100_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_7, data_out=>output_MAC_100_7);

	MAC_100_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_8, data_out=>output_MAC_100_8);

	MAC_100_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_9, data_out=>output_MAC_100_9);

	MAC_100_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_10, data_out=>output_MAC_100_10);

	MAC_100_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_11, data_out=>output_MAC_100_11);

	MAC_100_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_12, data_out=>output_MAC_100_12);

	MAC_100_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_13, data_out=>output_MAC_100_13);

	MAC_100_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_14, data_out=>output_MAC_100_14);

	MAC_100_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_15, data_out=>output_MAC_100_15);

	MAC_100_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_16, data_out=>output_MAC_100_16);

	MAC_100_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_17, data_out=>output_MAC_100_17);

	MAC_100_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_18, data_out=>output_MAC_100_18);

	MAC_100_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_19, data_out=>output_MAC_100_19);

	MAC_100_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_20, data_out=>output_MAC_100_20);

	MAC_100_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_21, data_out=>output_MAC_100_21);

	MAC_100_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_22, data_out=>output_MAC_100_22);

	MAC_100_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_23, data_out=>output_MAC_100_23);

	MAC_100_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_24, data_out=>output_MAC_100_24);

	MAC_100_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_25, data_out=>output_MAC_100_25);

	MAC_100_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_26, data_out=>output_MAC_100_26);

	MAC_100_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_27, data_out=>output_MAC_100_27);

	MAC_100_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_28, data_out=>output_MAC_100_28);

	MAC_100_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_29, data_out=>output_MAC_100_29);

	MAC_100_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_30, data_out=>output_MAC_100_30);

	MAC_100_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_100, data_in_B=>reg_input_col_31, data_out=>output_MAC_100_31);

	MAC_101_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_0, data_out=>output_MAC_101_0);

	MAC_101_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_1, data_out=>output_MAC_101_1);

	MAC_101_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_2, data_out=>output_MAC_101_2);

	MAC_101_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_3, data_out=>output_MAC_101_3);

	MAC_101_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_4, data_out=>output_MAC_101_4);

	MAC_101_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_5, data_out=>output_MAC_101_5);

	MAC_101_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_6, data_out=>output_MAC_101_6);

	MAC_101_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_7, data_out=>output_MAC_101_7);

	MAC_101_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_8, data_out=>output_MAC_101_8);

	MAC_101_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_9, data_out=>output_MAC_101_9);

	MAC_101_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_10, data_out=>output_MAC_101_10);

	MAC_101_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_11, data_out=>output_MAC_101_11);

	MAC_101_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_12, data_out=>output_MAC_101_12);

	MAC_101_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_13, data_out=>output_MAC_101_13);

	MAC_101_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_14, data_out=>output_MAC_101_14);

	MAC_101_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_15, data_out=>output_MAC_101_15);

	MAC_101_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_16, data_out=>output_MAC_101_16);

	MAC_101_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_17, data_out=>output_MAC_101_17);

	MAC_101_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_18, data_out=>output_MAC_101_18);

	MAC_101_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_19, data_out=>output_MAC_101_19);

	MAC_101_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_20, data_out=>output_MAC_101_20);

	MAC_101_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_21, data_out=>output_MAC_101_21);

	MAC_101_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_22, data_out=>output_MAC_101_22);

	MAC_101_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_23, data_out=>output_MAC_101_23);

	MAC_101_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_24, data_out=>output_MAC_101_24);

	MAC_101_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_25, data_out=>output_MAC_101_25);

	MAC_101_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_26, data_out=>output_MAC_101_26);

	MAC_101_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_27, data_out=>output_MAC_101_27);

	MAC_101_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_28, data_out=>output_MAC_101_28);

	MAC_101_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_29, data_out=>output_MAC_101_29);

	MAC_101_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_30, data_out=>output_MAC_101_30);

	MAC_101_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_101, data_in_B=>reg_input_col_31, data_out=>output_MAC_101_31);

	MAC_102_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_0, data_out=>output_MAC_102_0);

	MAC_102_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_1, data_out=>output_MAC_102_1);

	MAC_102_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_2, data_out=>output_MAC_102_2);

	MAC_102_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_3, data_out=>output_MAC_102_3);

	MAC_102_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_4, data_out=>output_MAC_102_4);

	MAC_102_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_5, data_out=>output_MAC_102_5);

	MAC_102_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_6, data_out=>output_MAC_102_6);

	MAC_102_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_7, data_out=>output_MAC_102_7);

	MAC_102_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_8, data_out=>output_MAC_102_8);

	MAC_102_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_9, data_out=>output_MAC_102_9);

	MAC_102_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_10, data_out=>output_MAC_102_10);

	MAC_102_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_11, data_out=>output_MAC_102_11);

	MAC_102_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_12, data_out=>output_MAC_102_12);

	MAC_102_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_13, data_out=>output_MAC_102_13);

	MAC_102_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_14, data_out=>output_MAC_102_14);

	MAC_102_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_15, data_out=>output_MAC_102_15);

	MAC_102_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_16, data_out=>output_MAC_102_16);

	MAC_102_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_17, data_out=>output_MAC_102_17);

	MAC_102_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_18, data_out=>output_MAC_102_18);

	MAC_102_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_19, data_out=>output_MAC_102_19);

	MAC_102_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_20, data_out=>output_MAC_102_20);

	MAC_102_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_21, data_out=>output_MAC_102_21);

	MAC_102_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_22, data_out=>output_MAC_102_22);

	MAC_102_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_23, data_out=>output_MAC_102_23);

	MAC_102_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_24, data_out=>output_MAC_102_24);

	MAC_102_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_25, data_out=>output_MAC_102_25);

	MAC_102_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_26, data_out=>output_MAC_102_26);

	MAC_102_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_27, data_out=>output_MAC_102_27);

	MAC_102_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_28, data_out=>output_MAC_102_28);

	MAC_102_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_29, data_out=>output_MAC_102_29);

	MAC_102_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_30, data_out=>output_MAC_102_30);

	MAC_102_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_102, data_in_B=>reg_input_col_31, data_out=>output_MAC_102_31);

	MAC_103_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_0, data_out=>output_MAC_103_0);

	MAC_103_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_1, data_out=>output_MAC_103_1);

	MAC_103_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_2, data_out=>output_MAC_103_2);

	MAC_103_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_3, data_out=>output_MAC_103_3);

	MAC_103_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_4, data_out=>output_MAC_103_4);

	MAC_103_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_5, data_out=>output_MAC_103_5);

	MAC_103_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_6, data_out=>output_MAC_103_6);

	MAC_103_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_7, data_out=>output_MAC_103_7);

	MAC_103_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_8, data_out=>output_MAC_103_8);

	MAC_103_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_9, data_out=>output_MAC_103_9);

	MAC_103_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_10, data_out=>output_MAC_103_10);

	MAC_103_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_11, data_out=>output_MAC_103_11);

	MAC_103_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_12, data_out=>output_MAC_103_12);

	MAC_103_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_13, data_out=>output_MAC_103_13);

	MAC_103_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_14, data_out=>output_MAC_103_14);

	MAC_103_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_15, data_out=>output_MAC_103_15);

	MAC_103_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_16, data_out=>output_MAC_103_16);

	MAC_103_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_17, data_out=>output_MAC_103_17);

	MAC_103_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_18, data_out=>output_MAC_103_18);

	MAC_103_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_19, data_out=>output_MAC_103_19);

	MAC_103_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_20, data_out=>output_MAC_103_20);

	MAC_103_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_21, data_out=>output_MAC_103_21);

	MAC_103_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_22, data_out=>output_MAC_103_22);

	MAC_103_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_23, data_out=>output_MAC_103_23);

	MAC_103_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_24, data_out=>output_MAC_103_24);

	MAC_103_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_25, data_out=>output_MAC_103_25);

	MAC_103_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_26, data_out=>output_MAC_103_26);

	MAC_103_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_27, data_out=>output_MAC_103_27);

	MAC_103_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_28, data_out=>output_MAC_103_28);

	MAC_103_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_29, data_out=>output_MAC_103_29);

	MAC_103_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_30, data_out=>output_MAC_103_30);

	MAC_103_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_103, data_in_B=>reg_input_col_31, data_out=>output_MAC_103_31);

	MAC_104_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_0, data_out=>output_MAC_104_0);

	MAC_104_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_1, data_out=>output_MAC_104_1);

	MAC_104_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_2, data_out=>output_MAC_104_2);

	MAC_104_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_3, data_out=>output_MAC_104_3);

	MAC_104_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_4, data_out=>output_MAC_104_4);

	MAC_104_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_5, data_out=>output_MAC_104_5);

	MAC_104_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_6, data_out=>output_MAC_104_6);

	MAC_104_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_7, data_out=>output_MAC_104_7);

	MAC_104_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_8, data_out=>output_MAC_104_8);

	MAC_104_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_9, data_out=>output_MAC_104_9);

	MAC_104_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_10, data_out=>output_MAC_104_10);

	MAC_104_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_11, data_out=>output_MAC_104_11);

	MAC_104_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_12, data_out=>output_MAC_104_12);

	MAC_104_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_13, data_out=>output_MAC_104_13);

	MAC_104_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_14, data_out=>output_MAC_104_14);

	MAC_104_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_15, data_out=>output_MAC_104_15);

	MAC_104_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_16, data_out=>output_MAC_104_16);

	MAC_104_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_17, data_out=>output_MAC_104_17);

	MAC_104_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_18, data_out=>output_MAC_104_18);

	MAC_104_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_19, data_out=>output_MAC_104_19);

	MAC_104_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_20, data_out=>output_MAC_104_20);

	MAC_104_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_21, data_out=>output_MAC_104_21);

	MAC_104_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_22, data_out=>output_MAC_104_22);

	MAC_104_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_23, data_out=>output_MAC_104_23);

	MAC_104_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_24, data_out=>output_MAC_104_24);

	MAC_104_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_25, data_out=>output_MAC_104_25);

	MAC_104_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_26, data_out=>output_MAC_104_26);

	MAC_104_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_27, data_out=>output_MAC_104_27);

	MAC_104_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_28, data_out=>output_MAC_104_28);

	MAC_104_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_29, data_out=>output_MAC_104_29);

	MAC_104_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_30, data_out=>output_MAC_104_30);

	MAC_104_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_104, data_in_B=>reg_input_col_31, data_out=>output_MAC_104_31);

	MAC_105_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_0, data_out=>output_MAC_105_0);

	MAC_105_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_1, data_out=>output_MAC_105_1);

	MAC_105_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_2, data_out=>output_MAC_105_2);

	MAC_105_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_3, data_out=>output_MAC_105_3);

	MAC_105_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_4, data_out=>output_MAC_105_4);

	MAC_105_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_5, data_out=>output_MAC_105_5);

	MAC_105_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_6, data_out=>output_MAC_105_6);

	MAC_105_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_7, data_out=>output_MAC_105_7);

	MAC_105_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_8, data_out=>output_MAC_105_8);

	MAC_105_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_9, data_out=>output_MAC_105_9);

	MAC_105_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_10, data_out=>output_MAC_105_10);

	MAC_105_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_11, data_out=>output_MAC_105_11);

	MAC_105_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_12, data_out=>output_MAC_105_12);

	MAC_105_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_13, data_out=>output_MAC_105_13);

	MAC_105_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_14, data_out=>output_MAC_105_14);

	MAC_105_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_15, data_out=>output_MAC_105_15);

	MAC_105_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_16, data_out=>output_MAC_105_16);

	MAC_105_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_17, data_out=>output_MAC_105_17);

	MAC_105_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_18, data_out=>output_MAC_105_18);

	MAC_105_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_19, data_out=>output_MAC_105_19);

	MAC_105_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_20, data_out=>output_MAC_105_20);

	MAC_105_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_21, data_out=>output_MAC_105_21);

	MAC_105_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_22, data_out=>output_MAC_105_22);

	MAC_105_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_23, data_out=>output_MAC_105_23);

	MAC_105_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_24, data_out=>output_MAC_105_24);

	MAC_105_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_25, data_out=>output_MAC_105_25);

	MAC_105_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_26, data_out=>output_MAC_105_26);

	MAC_105_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_27, data_out=>output_MAC_105_27);

	MAC_105_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_28, data_out=>output_MAC_105_28);

	MAC_105_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_29, data_out=>output_MAC_105_29);

	MAC_105_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_30, data_out=>output_MAC_105_30);

	MAC_105_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_105, data_in_B=>reg_input_col_31, data_out=>output_MAC_105_31);

	MAC_106_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_0, data_out=>output_MAC_106_0);

	MAC_106_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_1, data_out=>output_MAC_106_1);

	MAC_106_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_2, data_out=>output_MAC_106_2);

	MAC_106_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_3, data_out=>output_MAC_106_3);

	MAC_106_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_4, data_out=>output_MAC_106_4);

	MAC_106_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_5, data_out=>output_MAC_106_5);

	MAC_106_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_6, data_out=>output_MAC_106_6);

	MAC_106_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_7, data_out=>output_MAC_106_7);

	MAC_106_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_8, data_out=>output_MAC_106_8);

	MAC_106_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_9, data_out=>output_MAC_106_9);

	MAC_106_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_10, data_out=>output_MAC_106_10);

	MAC_106_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_11, data_out=>output_MAC_106_11);

	MAC_106_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_12, data_out=>output_MAC_106_12);

	MAC_106_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_13, data_out=>output_MAC_106_13);

	MAC_106_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_14, data_out=>output_MAC_106_14);

	MAC_106_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_15, data_out=>output_MAC_106_15);

	MAC_106_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_16, data_out=>output_MAC_106_16);

	MAC_106_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_17, data_out=>output_MAC_106_17);

	MAC_106_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_18, data_out=>output_MAC_106_18);

	MAC_106_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_19, data_out=>output_MAC_106_19);

	MAC_106_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_20, data_out=>output_MAC_106_20);

	MAC_106_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_21, data_out=>output_MAC_106_21);

	MAC_106_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_22, data_out=>output_MAC_106_22);

	MAC_106_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_23, data_out=>output_MAC_106_23);

	MAC_106_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_24, data_out=>output_MAC_106_24);

	MAC_106_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_25, data_out=>output_MAC_106_25);

	MAC_106_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_26, data_out=>output_MAC_106_26);

	MAC_106_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_27, data_out=>output_MAC_106_27);

	MAC_106_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_28, data_out=>output_MAC_106_28);

	MAC_106_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_29, data_out=>output_MAC_106_29);

	MAC_106_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_30, data_out=>output_MAC_106_30);

	MAC_106_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_106, data_in_B=>reg_input_col_31, data_out=>output_MAC_106_31);

	MAC_107_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_0, data_out=>output_MAC_107_0);

	MAC_107_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_1, data_out=>output_MAC_107_1);

	MAC_107_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_2, data_out=>output_MAC_107_2);

	MAC_107_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_3, data_out=>output_MAC_107_3);

	MAC_107_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_4, data_out=>output_MAC_107_4);

	MAC_107_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_5, data_out=>output_MAC_107_5);

	MAC_107_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_6, data_out=>output_MAC_107_6);

	MAC_107_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_7, data_out=>output_MAC_107_7);

	MAC_107_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_8, data_out=>output_MAC_107_8);

	MAC_107_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_9, data_out=>output_MAC_107_9);

	MAC_107_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_10, data_out=>output_MAC_107_10);

	MAC_107_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_11, data_out=>output_MAC_107_11);

	MAC_107_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_12, data_out=>output_MAC_107_12);

	MAC_107_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_13, data_out=>output_MAC_107_13);

	MAC_107_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_14, data_out=>output_MAC_107_14);

	MAC_107_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_15, data_out=>output_MAC_107_15);

	MAC_107_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_16, data_out=>output_MAC_107_16);

	MAC_107_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_17, data_out=>output_MAC_107_17);

	MAC_107_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_18, data_out=>output_MAC_107_18);

	MAC_107_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_19, data_out=>output_MAC_107_19);

	MAC_107_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_20, data_out=>output_MAC_107_20);

	MAC_107_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_21, data_out=>output_MAC_107_21);

	MAC_107_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_22, data_out=>output_MAC_107_22);

	MAC_107_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_23, data_out=>output_MAC_107_23);

	MAC_107_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_24, data_out=>output_MAC_107_24);

	MAC_107_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_25, data_out=>output_MAC_107_25);

	MAC_107_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_26, data_out=>output_MAC_107_26);

	MAC_107_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_27, data_out=>output_MAC_107_27);

	MAC_107_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_28, data_out=>output_MAC_107_28);

	MAC_107_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_29, data_out=>output_MAC_107_29);

	MAC_107_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_30, data_out=>output_MAC_107_30);

	MAC_107_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_107, data_in_B=>reg_input_col_31, data_out=>output_MAC_107_31);

	MAC_108_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_0, data_out=>output_MAC_108_0);

	MAC_108_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_1, data_out=>output_MAC_108_1);

	MAC_108_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_2, data_out=>output_MAC_108_2);

	MAC_108_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_3, data_out=>output_MAC_108_3);

	MAC_108_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_4, data_out=>output_MAC_108_4);

	MAC_108_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_5, data_out=>output_MAC_108_5);

	MAC_108_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_6, data_out=>output_MAC_108_6);

	MAC_108_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_7, data_out=>output_MAC_108_7);

	MAC_108_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_8, data_out=>output_MAC_108_8);

	MAC_108_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_9, data_out=>output_MAC_108_9);

	MAC_108_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_10, data_out=>output_MAC_108_10);

	MAC_108_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_11, data_out=>output_MAC_108_11);

	MAC_108_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_12, data_out=>output_MAC_108_12);

	MAC_108_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_13, data_out=>output_MAC_108_13);

	MAC_108_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_14, data_out=>output_MAC_108_14);

	MAC_108_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_15, data_out=>output_MAC_108_15);

	MAC_108_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_16, data_out=>output_MAC_108_16);

	MAC_108_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_17, data_out=>output_MAC_108_17);

	MAC_108_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_18, data_out=>output_MAC_108_18);

	MAC_108_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_19, data_out=>output_MAC_108_19);

	MAC_108_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_20, data_out=>output_MAC_108_20);

	MAC_108_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_21, data_out=>output_MAC_108_21);

	MAC_108_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_22, data_out=>output_MAC_108_22);

	MAC_108_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_23, data_out=>output_MAC_108_23);

	MAC_108_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_24, data_out=>output_MAC_108_24);

	MAC_108_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_25, data_out=>output_MAC_108_25);

	MAC_108_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_26, data_out=>output_MAC_108_26);

	MAC_108_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_27, data_out=>output_MAC_108_27);

	MAC_108_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_28, data_out=>output_MAC_108_28);

	MAC_108_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_29, data_out=>output_MAC_108_29);

	MAC_108_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_30, data_out=>output_MAC_108_30);

	MAC_108_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_108, data_in_B=>reg_input_col_31, data_out=>output_MAC_108_31);

	MAC_109_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_0, data_out=>output_MAC_109_0);

	MAC_109_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_1, data_out=>output_MAC_109_1);

	MAC_109_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_2, data_out=>output_MAC_109_2);

	MAC_109_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_3, data_out=>output_MAC_109_3);

	MAC_109_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_4, data_out=>output_MAC_109_4);

	MAC_109_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_5, data_out=>output_MAC_109_5);

	MAC_109_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_6, data_out=>output_MAC_109_6);

	MAC_109_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_7, data_out=>output_MAC_109_7);

	MAC_109_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_8, data_out=>output_MAC_109_8);

	MAC_109_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_9, data_out=>output_MAC_109_9);

	MAC_109_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_10, data_out=>output_MAC_109_10);

	MAC_109_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_11, data_out=>output_MAC_109_11);

	MAC_109_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_12, data_out=>output_MAC_109_12);

	MAC_109_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_13, data_out=>output_MAC_109_13);

	MAC_109_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_14, data_out=>output_MAC_109_14);

	MAC_109_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_15, data_out=>output_MAC_109_15);

	MAC_109_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_16, data_out=>output_MAC_109_16);

	MAC_109_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_17, data_out=>output_MAC_109_17);

	MAC_109_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_18, data_out=>output_MAC_109_18);

	MAC_109_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_19, data_out=>output_MAC_109_19);

	MAC_109_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_20, data_out=>output_MAC_109_20);

	MAC_109_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_21, data_out=>output_MAC_109_21);

	MAC_109_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_22, data_out=>output_MAC_109_22);

	MAC_109_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_23, data_out=>output_MAC_109_23);

	MAC_109_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_24, data_out=>output_MAC_109_24);

	MAC_109_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_25, data_out=>output_MAC_109_25);

	MAC_109_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_26, data_out=>output_MAC_109_26);

	MAC_109_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_27, data_out=>output_MAC_109_27);

	MAC_109_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_28, data_out=>output_MAC_109_28);

	MAC_109_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_29, data_out=>output_MAC_109_29);

	MAC_109_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_30, data_out=>output_MAC_109_30);

	MAC_109_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_109, data_in_B=>reg_input_col_31, data_out=>output_MAC_109_31);

	MAC_110_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_0, data_out=>output_MAC_110_0);

	MAC_110_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_1, data_out=>output_MAC_110_1);

	MAC_110_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_2, data_out=>output_MAC_110_2);

	MAC_110_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_3, data_out=>output_MAC_110_3);

	MAC_110_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_4, data_out=>output_MAC_110_4);

	MAC_110_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_5, data_out=>output_MAC_110_5);

	MAC_110_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_6, data_out=>output_MAC_110_6);

	MAC_110_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_7, data_out=>output_MAC_110_7);

	MAC_110_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_8, data_out=>output_MAC_110_8);

	MAC_110_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_9, data_out=>output_MAC_110_9);

	MAC_110_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_10, data_out=>output_MAC_110_10);

	MAC_110_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_11, data_out=>output_MAC_110_11);

	MAC_110_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_12, data_out=>output_MAC_110_12);

	MAC_110_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_13, data_out=>output_MAC_110_13);

	MAC_110_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_14, data_out=>output_MAC_110_14);

	MAC_110_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_15, data_out=>output_MAC_110_15);

	MAC_110_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_16, data_out=>output_MAC_110_16);

	MAC_110_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_17, data_out=>output_MAC_110_17);

	MAC_110_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_18, data_out=>output_MAC_110_18);

	MAC_110_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_19, data_out=>output_MAC_110_19);

	MAC_110_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_20, data_out=>output_MAC_110_20);

	MAC_110_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_21, data_out=>output_MAC_110_21);

	MAC_110_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_22, data_out=>output_MAC_110_22);

	MAC_110_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_23, data_out=>output_MAC_110_23);

	MAC_110_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_24, data_out=>output_MAC_110_24);

	MAC_110_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_25, data_out=>output_MAC_110_25);

	MAC_110_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_26, data_out=>output_MAC_110_26);

	MAC_110_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_27, data_out=>output_MAC_110_27);

	MAC_110_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_28, data_out=>output_MAC_110_28);

	MAC_110_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_29, data_out=>output_MAC_110_29);

	MAC_110_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_30, data_out=>output_MAC_110_30);

	MAC_110_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_110, data_in_B=>reg_input_col_31, data_out=>output_MAC_110_31);

	MAC_111_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_0, data_out=>output_MAC_111_0);

	MAC_111_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_1, data_out=>output_MAC_111_1);

	MAC_111_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_2, data_out=>output_MAC_111_2);

	MAC_111_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_3, data_out=>output_MAC_111_3);

	MAC_111_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_4, data_out=>output_MAC_111_4);

	MAC_111_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_5, data_out=>output_MAC_111_5);

	MAC_111_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_6, data_out=>output_MAC_111_6);

	MAC_111_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_7, data_out=>output_MAC_111_7);

	MAC_111_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_8, data_out=>output_MAC_111_8);

	MAC_111_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_9, data_out=>output_MAC_111_9);

	MAC_111_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_10, data_out=>output_MAC_111_10);

	MAC_111_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_11, data_out=>output_MAC_111_11);

	MAC_111_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_12, data_out=>output_MAC_111_12);

	MAC_111_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_13, data_out=>output_MAC_111_13);

	MAC_111_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_14, data_out=>output_MAC_111_14);

	MAC_111_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_15, data_out=>output_MAC_111_15);

	MAC_111_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_16, data_out=>output_MAC_111_16);

	MAC_111_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_17, data_out=>output_MAC_111_17);

	MAC_111_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_18, data_out=>output_MAC_111_18);

	MAC_111_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_19, data_out=>output_MAC_111_19);

	MAC_111_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_20, data_out=>output_MAC_111_20);

	MAC_111_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_21, data_out=>output_MAC_111_21);

	MAC_111_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_22, data_out=>output_MAC_111_22);

	MAC_111_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_23, data_out=>output_MAC_111_23);

	MAC_111_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_24, data_out=>output_MAC_111_24);

	MAC_111_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_25, data_out=>output_MAC_111_25);

	MAC_111_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_26, data_out=>output_MAC_111_26);

	MAC_111_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_27, data_out=>output_MAC_111_27);

	MAC_111_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_28, data_out=>output_MAC_111_28);

	MAC_111_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_29, data_out=>output_MAC_111_29);

	MAC_111_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_30, data_out=>output_MAC_111_30);

	MAC_111_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_111, data_in_B=>reg_input_col_31, data_out=>output_MAC_111_31);

	MAC_112_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_0, data_out=>output_MAC_112_0);

	MAC_112_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_1, data_out=>output_MAC_112_1);

	MAC_112_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_2, data_out=>output_MAC_112_2);

	MAC_112_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_3, data_out=>output_MAC_112_3);

	MAC_112_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_4, data_out=>output_MAC_112_4);

	MAC_112_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_5, data_out=>output_MAC_112_5);

	MAC_112_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_6, data_out=>output_MAC_112_6);

	MAC_112_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_7, data_out=>output_MAC_112_7);

	MAC_112_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_8, data_out=>output_MAC_112_8);

	MAC_112_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_9, data_out=>output_MAC_112_9);

	MAC_112_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_10, data_out=>output_MAC_112_10);

	MAC_112_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_11, data_out=>output_MAC_112_11);

	MAC_112_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_12, data_out=>output_MAC_112_12);

	MAC_112_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_13, data_out=>output_MAC_112_13);

	MAC_112_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_14, data_out=>output_MAC_112_14);

	MAC_112_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_15, data_out=>output_MAC_112_15);

	MAC_112_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_16, data_out=>output_MAC_112_16);

	MAC_112_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_17, data_out=>output_MAC_112_17);

	MAC_112_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_18, data_out=>output_MAC_112_18);

	MAC_112_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_19, data_out=>output_MAC_112_19);

	MAC_112_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_20, data_out=>output_MAC_112_20);

	MAC_112_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_21, data_out=>output_MAC_112_21);

	MAC_112_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_22, data_out=>output_MAC_112_22);

	MAC_112_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_23, data_out=>output_MAC_112_23);

	MAC_112_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_24, data_out=>output_MAC_112_24);

	MAC_112_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_25, data_out=>output_MAC_112_25);

	MAC_112_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_26, data_out=>output_MAC_112_26);

	MAC_112_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_27, data_out=>output_MAC_112_27);

	MAC_112_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_28, data_out=>output_MAC_112_28);

	MAC_112_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_29, data_out=>output_MAC_112_29);

	MAC_112_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_30, data_out=>output_MAC_112_30);

	MAC_112_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_112, data_in_B=>reg_input_col_31, data_out=>output_MAC_112_31);

	MAC_113_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_0, data_out=>output_MAC_113_0);

	MAC_113_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_1, data_out=>output_MAC_113_1);

	MAC_113_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_2, data_out=>output_MAC_113_2);

	MAC_113_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_3, data_out=>output_MAC_113_3);

	MAC_113_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_4, data_out=>output_MAC_113_4);

	MAC_113_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_5, data_out=>output_MAC_113_5);

	MAC_113_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_6, data_out=>output_MAC_113_6);

	MAC_113_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_7, data_out=>output_MAC_113_7);

	MAC_113_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_8, data_out=>output_MAC_113_8);

	MAC_113_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_9, data_out=>output_MAC_113_9);

	MAC_113_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_10, data_out=>output_MAC_113_10);

	MAC_113_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_11, data_out=>output_MAC_113_11);

	MAC_113_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_12, data_out=>output_MAC_113_12);

	MAC_113_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_13, data_out=>output_MAC_113_13);

	MAC_113_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_14, data_out=>output_MAC_113_14);

	MAC_113_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_15, data_out=>output_MAC_113_15);

	MAC_113_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_16, data_out=>output_MAC_113_16);

	MAC_113_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_17, data_out=>output_MAC_113_17);

	MAC_113_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_18, data_out=>output_MAC_113_18);

	MAC_113_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_19, data_out=>output_MAC_113_19);

	MAC_113_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_20, data_out=>output_MAC_113_20);

	MAC_113_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_21, data_out=>output_MAC_113_21);

	MAC_113_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_22, data_out=>output_MAC_113_22);

	MAC_113_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_23, data_out=>output_MAC_113_23);

	MAC_113_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_24, data_out=>output_MAC_113_24);

	MAC_113_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_25, data_out=>output_MAC_113_25);

	MAC_113_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_26, data_out=>output_MAC_113_26);

	MAC_113_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_27, data_out=>output_MAC_113_27);

	MAC_113_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_28, data_out=>output_MAC_113_28);

	MAC_113_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_29, data_out=>output_MAC_113_29);

	MAC_113_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_30, data_out=>output_MAC_113_30);

	MAC_113_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_113, data_in_B=>reg_input_col_31, data_out=>output_MAC_113_31);

	MAC_114_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_0, data_out=>output_MAC_114_0);

	MAC_114_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_1, data_out=>output_MAC_114_1);

	MAC_114_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_2, data_out=>output_MAC_114_2);

	MAC_114_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_3, data_out=>output_MAC_114_3);

	MAC_114_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_4, data_out=>output_MAC_114_4);

	MAC_114_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_5, data_out=>output_MAC_114_5);

	MAC_114_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_6, data_out=>output_MAC_114_6);

	MAC_114_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_7, data_out=>output_MAC_114_7);

	MAC_114_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_8, data_out=>output_MAC_114_8);

	MAC_114_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_9, data_out=>output_MAC_114_9);

	MAC_114_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_10, data_out=>output_MAC_114_10);

	MAC_114_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_11, data_out=>output_MAC_114_11);

	MAC_114_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_12, data_out=>output_MAC_114_12);

	MAC_114_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_13, data_out=>output_MAC_114_13);

	MAC_114_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_14, data_out=>output_MAC_114_14);

	MAC_114_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_15, data_out=>output_MAC_114_15);

	MAC_114_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_16, data_out=>output_MAC_114_16);

	MAC_114_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_17, data_out=>output_MAC_114_17);

	MAC_114_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_18, data_out=>output_MAC_114_18);

	MAC_114_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_19, data_out=>output_MAC_114_19);

	MAC_114_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_20, data_out=>output_MAC_114_20);

	MAC_114_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_21, data_out=>output_MAC_114_21);

	MAC_114_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_22, data_out=>output_MAC_114_22);

	MAC_114_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_23, data_out=>output_MAC_114_23);

	MAC_114_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_24, data_out=>output_MAC_114_24);

	MAC_114_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_25, data_out=>output_MAC_114_25);

	MAC_114_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_26, data_out=>output_MAC_114_26);

	MAC_114_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_27, data_out=>output_MAC_114_27);

	MAC_114_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_28, data_out=>output_MAC_114_28);

	MAC_114_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_29, data_out=>output_MAC_114_29);

	MAC_114_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_30, data_out=>output_MAC_114_30);

	MAC_114_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_114, data_in_B=>reg_input_col_31, data_out=>output_MAC_114_31);

	MAC_115_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_0, data_out=>output_MAC_115_0);

	MAC_115_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_1, data_out=>output_MAC_115_1);

	MAC_115_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_2, data_out=>output_MAC_115_2);

	MAC_115_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_3, data_out=>output_MAC_115_3);

	MAC_115_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_4, data_out=>output_MAC_115_4);

	MAC_115_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_5, data_out=>output_MAC_115_5);

	MAC_115_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_6, data_out=>output_MAC_115_6);

	MAC_115_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_7, data_out=>output_MAC_115_7);

	MAC_115_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_8, data_out=>output_MAC_115_8);

	MAC_115_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_9, data_out=>output_MAC_115_9);

	MAC_115_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_10, data_out=>output_MAC_115_10);

	MAC_115_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_11, data_out=>output_MAC_115_11);

	MAC_115_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_12, data_out=>output_MAC_115_12);

	MAC_115_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_13, data_out=>output_MAC_115_13);

	MAC_115_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_14, data_out=>output_MAC_115_14);

	MAC_115_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_15, data_out=>output_MAC_115_15);

	MAC_115_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_16, data_out=>output_MAC_115_16);

	MAC_115_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_17, data_out=>output_MAC_115_17);

	MAC_115_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_18, data_out=>output_MAC_115_18);

	MAC_115_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_19, data_out=>output_MAC_115_19);

	MAC_115_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_20, data_out=>output_MAC_115_20);

	MAC_115_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_21, data_out=>output_MAC_115_21);

	MAC_115_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_22, data_out=>output_MAC_115_22);

	MAC_115_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_23, data_out=>output_MAC_115_23);

	MAC_115_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_24, data_out=>output_MAC_115_24);

	MAC_115_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_25, data_out=>output_MAC_115_25);

	MAC_115_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_26, data_out=>output_MAC_115_26);

	MAC_115_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_27, data_out=>output_MAC_115_27);

	MAC_115_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_28, data_out=>output_MAC_115_28);

	MAC_115_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_29, data_out=>output_MAC_115_29);

	MAC_115_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_30, data_out=>output_MAC_115_30);

	MAC_115_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_115, data_in_B=>reg_input_col_31, data_out=>output_MAC_115_31);

	MAC_116_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_0, data_out=>output_MAC_116_0);

	MAC_116_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_1, data_out=>output_MAC_116_1);

	MAC_116_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_2, data_out=>output_MAC_116_2);

	MAC_116_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_3, data_out=>output_MAC_116_3);

	MAC_116_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_4, data_out=>output_MAC_116_4);

	MAC_116_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_5, data_out=>output_MAC_116_5);

	MAC_116_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_6, data_out=>output_MAC_116_6);

	MAC_116_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_7, data_out=>output_MAC_116_7);

	MAC_116_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_8, data_out=>output_MAC_116_8);

	MAC_116_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_9, data_out=>output_MAC_116_9);

	MAC_116_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_10, data_out=>output_MAC_116_10);

	MAC_116_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_11, data_out=>output_MAC_116_11);

	MAC_116_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_12, data_out=>output_MAC_116_12);

	MAC_116_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_13, data_out=>output_MAC_116_13);

	MAC_116_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_14, data_out=>output_MAC_116_14);

	MAC_116_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_15, data_out=>output_MAC_116_15);

	MAC_116_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_16, data_out=>output_MAC_116_16);

	MAC_116_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_17, data_out=>output_MAC_116_17);

	MAC_116_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_18, data_out=>output_MAC_116_18);

	MAC_116_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_19, data_out=>output_MAC_116_19);

	MAC_116_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_20, data_out=>output_MAC_116_20);

	MAC_116_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_21, data_out=>output_MAC_116_21);

	MAC_116_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_22, data_out=>output_MAC_116_22);

	MAC_116_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_23, data_out=>output_MAC_116_23);

	MAC_116_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_24, data_out=>output_MAC_116_24);

	MAC_116_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_25, data_out=>output_MAC_116_25);

	MAC_116_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_26, data_out=>output_MAC_116_26);

	MAC_116_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_27, data_out=>output_MAC_116_27);

	MAC_116_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_28, data_out=>output_MAC_116_28);

	MAC_116_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_29, data_out=>output_MAC_116_29);

	MAC_116_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_30, data_out=>output_MAC_116_30);

	MAC_116_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_116, data_in_B=>reg_input_col_31, data_out=>output_MAC_116_31);

	MAC_117_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_0, data_out=>output_MAC_117_0);

	MAC_117_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_1, data_out=>output_MAC_117_1);

	MAC_117_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_2, data_out=>output_MAC_117_2);

	MAC_117_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_3, data_out=>output_MAC_117_3);

	MAC_117_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_4, data_out=>output_MAC_117_4);

	MAC_117_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_5, data_out=>output_MAC_117_5);

	MAC_117_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_6, data_out=>output_MAC_117_6);

	MAC_117_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_7, data_out=>output_MAC_117_7);

	MAC_117_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_8, data_out=>output_MAC_117_8);

	MAC_117_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_9, data_out=>output_MAC_117_9);

	MAC_117_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_10, data_out=>output_MAC_117_10);

	MAC_117_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_11, data_out=>output_MAC_117_11);

	MAC_117_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_12, data_out=>output_MAC_117_12);

	MAC_117_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_13, data_out=>output_MAC_117_13);

	MAC_117_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_14, data_out=>output_MAC_117_14);

	MAC_117_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_15, data_out=>output_MAC_117_15);

	MAC_117_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_16, data_out=>output_MAC_117_16);

	MAC_117_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_17, data_out=>output_MAC_117_17);

	MAC_117_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_18, data_out=>output_MAC_117_18);

	MAC_117_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_19, data_out=>output_MAC_117_19);

	MAC_117_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_20, data_out=>output_MAC_117_20);

	MAC_117_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_21, data_out=>output_MAC_117_21);

	MAC_117_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_22, data_out=>output_MAC_117_22);

	MAC_117_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_23, data_out=>output_MAC_117_23);

	MAC_117_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_24, data_out=>output_MAC_117_24);

	MAC_117_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_25, data_out=>output_MAC_117_25);

	MAC_117_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_26, data_out=>output_MAC_117_26);

	MAC_117_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_27, data_out=>output_MAC_117_27);

	MAC_117_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_28, data_out=>output_MAC_117_28);

	MAC_117_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_29, data_out=>output_MAC_117_29);

	MAC_117_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_30, data_out=>output_MAC_117_30);

	MAC_117_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_117, data_in_B=>reg_input_col_31, data_out=>output_MAC_117_31);

	MAC_118_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_0, data_out=>output_MAC_118_0);

	MAC_118_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_1, data_out=>output_MAC_118_1);

	MAC_118_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_2, data_out=>output_MAC_118_2);

	MAC_118_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_3, data_out=>output_MAC_118_3);

	MAC_118_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_4, data_out=>output_MAC_118_4);

	MAC_118_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_5, data_out=>output_MAC_118_5);

	MAC_118_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_6, data_out=>output_MAC_118_6);

	MAC_118_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_7, data_out=>output_MAC_118_7);

	MAC_118_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_8, data_out=>output_MAC_118_8);

	MAC_118_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_9, data_out=>output_MAC_118_9);

	MAC_118_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_10, data_out=>output_MAC_118_10);

	MAC_118_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_11, data_out=>output_MAC_118_11);

	MAC_118_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_12, data_out=>output_MAC_118_12);

	MAC_118_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_13, data_out=>output_MAC_118_13);

	MAC_118_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_14, data_out=>output_MAC_118_14);

	MAC_118_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_15, data_out=>output_MAC_118_15);

	MAC_118_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_16, data_out=>output_MAC_118_16);

	MAC_118_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_17, data_out=>output_MAC_118_17);

	MAC_118_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_18, data_out=>output_MAC_118_18);

	MAC_118_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_19, data_out=>output_MAC_118_19);

	MAC_118_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_20, data_out=>output_MAC_118_20);

	MAC_118_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_21, data_out=>output_MAC_118_21);

	MAC_118_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_22, data_out=>output_MAC_118_22);

	MAC_118_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_23, data_out=>output_MAC_118_23);

	MAC_118_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_24, data_out=>output_MAC_118_24);

	MAC_118_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_25, data_out=>output_MAC_118_25);

	MAC_118_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_26, data_out=>output_MAC_118_26);

	MAC_118_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_27, data_out=>output_MAC_118_27);

	MAC_118_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_28, data_out=>output_MAC_118_28);

	MAC_118_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_29, data_out=>output_MAC_118_29);

	MAC_118_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_30, data_out=>output_MAC_118_30);

	MAC_118_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_118, data_in_B=>reg_input_col_31, data_out=>output_MAC_118_31);

	MAC_119_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_0, data_out=>output_MAC_119_0);

	MAC_119_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_1, data_out=>output_MAC_119_1);

	MAC_119_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_2, data_out=>output_MAC_119_2);

	MAC_119_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_3, data_out=>output_MAC_119_3);

	MAC_119_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_4, data_out=>output_MAC_119_4);

	MAC_119_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_5, data_out=>output_MAC_119_5);

	MAC_119_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_6, data_out=>output_MAC_119_6);

	MAC_119_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_7, data_out=>output_MAC_119_7);

	MAC_119_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_8, data_out=>output_MAC_119_8);

	MAC_119_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_9, data_out=>output_MAC_119_9);

	MAC_119_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_10, data_out=>output_MAC_119_10);

	MAC_119_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_11, data_out=>output_MAC_119_11);

	MAC_119_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_12, data_out=>output_MAC_119_12);

	MAC_119_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_13, data_out=>output_MAC_119_13);

	MAC_119_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_14, data_out=>output_MAC_119_14);

	MAC_119_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_15, data_out=>output_MAC_119_15);

	MAC_119_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_16, data_out=>output_MAC_119_16);

	MAC_119_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_17, data_out=>output_MAC_119_17);

	MAC_119_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_18, data_out=>output_MAC_119_18);

	MAC_119_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_19, data_out=>output_MAC_119_19);

	MAC_119_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_20, data_out=>output_MAC_119_20);

	MAC_119_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_21, data_out=>output_MAC_119_21);

	MAC_119_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_22, data_out=>output_MAC_119_22);

	MAC_119_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_23, data_out=>output_MAC_119_23);

	MAC_119_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_24, data_out=>output_MAC_119_24);

	MAC_119_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_25, data_out=>output_MAC_119_25);

	MAC_119_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_26, data_out=>output_MAC_119_26);

	MAC_119_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_27, data_out=>output_MAC_119_27);

	MAC_119_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_28, data_out=>output_MAC_119_28);

	MAC_119_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_29, data_out=>output_MAC_119_29);

	MAC_119_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_30, data_out=>output_MAC_119_30);

	MAC_119_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_119, data_in_B=>reg_input_col_31, data_out=>output_MAC_119_31);

	MAC_120_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_0, data_out=>output_MAC_120_0);

	MAC_120_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_1, data_out=>output_MAC_120_1);

	MAC_120_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_2, data_out=>output_MAC_120_2);

	MAC_120_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_3, data_out=>output_MAC_120_3);

	MAC_120_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_4, data_out=>output_MAC_120_4);

	MAC_120_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_5, data_out=>output_MAC_120_5);

	MAC_120_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_6, data_out=>output_MAC_120_6);

	MAC_120_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_7, data_out=>output_MAC_120_7);

	MAC_120_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_8, data_out=>output_MAC_120_8);

	MAC_120_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_9, data_out=>output_MAC_120_9);

	MAC_120_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_10, data_out=>output_MAC_120_10);

	MAC_120_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_11, data_out=>output_MAC_120_11);

	MAC_120_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_12, data_out=>output_MAC_120_12);

	MAC_120_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_13, data_out=>output_MAC_120_13);

	MAC_120_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_14, data_out=>output_MAC_120_14);

	MAC_120_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_15, data_out=>output_MAC_120_15);

	MAC_120_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_16, data_out=>output_MAC_120_16);

	MAC_120_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_17, data_out=>output_MAC_120_17);

	MAC_120_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_18, data_out=>output_MAC_120_18);

	MAC_120_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_19, data_out=>output_MAC_120_19);

	MAC_120_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_20, data_out=>output_MAC_120_20);

	MAC_120_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_21, data_out=>output_MAC_120_21);

	MAC_120_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_22, data_out=>output_MAC_120_22);

	MAC_120_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_23, data_out=>output_MAC_120_23);

	MAC_120_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_24, data_out=>output_MAC_120_24);

	MAC_120_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_25, data_out=>output_MAC_120_25);

	MAC_120_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_26, data_out=>output_MAC_120_26);

	MAC_120_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_27, data_out=>output_MAC_120_27);

	MAC_120_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_28, data_out=>output_MAC_120_28);

	MAC_120_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_29, data_out=>output_MAC_120_29);

	MAC_120_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_30, data_out=>output_MAC_120_30);

	MAC_120_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_120, data_in_B=>reg_input_col_31, data_out=>output_MAC_120_31);

	MAC_121_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_0, data_out=>output_MAC_121_0);

	MAC_121_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_1, data_out=>output_MAC_121_1);

	MAC_121_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_2, data_out=>output_MAC_121_2);

	MAC_121_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_3, data_out=>output_MAC_121_3);

	MAC_121_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_4, data_out=>output_MAC_121_4);

	MAC_121_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_5, data_out=>output_MAC_121_5);

	MAC_121_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_6, data_out=>output_MAC_121_6);

	MAC_121_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_7, data_out=>output_MAC_121_7);

	MAC_121_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_8, data_out=>output_MAC_121_8);

	MAC_121_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_9, data_out=>output_MAC_121_9);

	MAC_121_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_10, data_out=>output_MAC_121_10);

	MAC_121_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_11, data_out=>output_MAC_121_11);

	MAC_121_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_12, data_out=>output_MAC_121_12);

	MAC_121_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_13, data_out=>output_MAC_121_13);

	MAC_121_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_14, data_out=>output_MAC_121_14);

	MAC_121_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_15, data_out=>output_MAC_121_15);

	MAC_121_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_16, data_out=>output_MAC_121_16);

	MAC_121_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_17, data_out=>output_MAC_121_17);

	MAC_121_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_18, data_out=>output_MAC_121_18);

	MAC_121_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_19, data_out=>output_MAC_121_19);

	MAC_121_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_20, data_out=>output_MAC_121_20);

	MAC_121_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_21, data_out=>output_MAC_121_21);

	MAC_121_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_22, data_out=>output_MAC_121_22);

	MAC_121_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_23, data_out=>output_MAC_121_23);

	MAC_121_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_24, data_out=>output_MAC_121_24);

	MAC_121_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_25, data_out=>output_MAC_121_25);

	MAC_121_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_26, data_out=>output_MAC_121_26);

	MAC_121_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_27, data_out=>output_MAC_121_27);

	MAC_121_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_28, data_out=>output_MAC_121_28);

	MAC_121_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_29, data_out=>output_MAC_121_29);

	MAC_121_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_30, data_out=>output_MAC_121_30);

	MAC_121_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_121, data_in_B=>reg_input_col_31, data_out=>output_MAC_121_31);

	MAC_122_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_0, data_out=>output_MAC_122_0);

	MAC_122_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_1, data_out=>output_MAC_122_1);

	MAC_122_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_2, data_out=>output_MAC_122_2);

	MAC_122_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_3, data_out=>output_MAC_122_3);

	MAC_122_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_4, data_out=>output_MAC_122_4);

	MAC_122_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_5, data_out=>output_MAC_122_5);

	MAC_122_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_6, data_out=>output_MAC_122_6);

	MAC_122_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_7, data_out=>output_MAC_122_7);

	MAC_122_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_8, data_out=>output_MAC_122_8);

	MAC_122_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_9, data_out=>output_MAC_122_9);

	MAC_122_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_10, data_out=>output_MAC_122_10);

	MAC_122_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_11, data_out=>output_MAC_122_11);

	MAC_122_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_12, data_out=>output_MAC_122_12);

	MAC_122_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_13, data_out=>output_MAC_122_13);

	MAC_122_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_14, data_out=>output_MAC_122_14);

	MAC_122_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_15, data_out=>output_MAC_122_15);

	MAC_122_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_16, data_out=>output_MAC_122_16);

	MAC_122_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_17, data_out=>output_MAC_122_17);

	MAC_122_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_18, data_out=>output_MAC_122_18);

	MAC_122_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_19, data_out=>output_MAC_122_19);

	MAC_122_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_20, data_out=>output_MAC_122_20);

	MAC_122_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_21, data_out=>output_MAC_122_21);

	MAC_122_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_22, data_out=>output_MAC_122_22);

	MAC_122_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_23, data_out=>output_MAC_122_23);

	MAC_122_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_24, data_out=>output_MAC_122_24);

	MAC_122_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_25, data_out=>output_MAC_122_25);

	MAC_122_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_26, data_out=>output_MAC_122_26);

	MAC_122_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_27, data_out=>output_MAC_122_27);

	MAC_122_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_28, data_out=>output_MAC_122_28);

	MAC_122_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_29, data_out=>output_MAC_122_29);

	MAC_122_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_30, data_out=>output_MAC_122_30);

	MAC_122_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_122, data_in_B=>reg_input_col_31, data_out=>output_MAC_122_31);

	MAC_123_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_0, data_out=>output_MAC_123_0);

	MAC_123_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_1, data_out=>output_MAC_123_1);

	MAC_123_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_2, data_out=>output_MAC_123_2);

	MAC_123_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_3, data_out=>output_MAC_123_3);

	MAC_123_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_4, data_out=>output_MAC_123_4);

	MAC_123_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_5, data_out=>output_MAC_123_5);

	MAC_123_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_6, data_out=>output_MAC_123_6);

	MAC_123_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_7, data_out=>output_MAC_123_7);

	MAC_123_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_8, data_out=>output_MAC_123_8);

	MAC_123_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_9, data_out=>output_MAC_123_9);

	MAC_123_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_10, data_out=>output_MAC_123_10);

	MAC_123_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_11, data_out=>output_MAC_123_11);

	MAC_123_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_12, data_out=>output_MAC_123_12);

	MAC_123_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_13, data_out=>output_MAC_123_13);

	MAC_123_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_14, data_out=>output_MAC_123_14);

	MAC_123_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_15, data_out=>output_MAC_123_15);

	MAC_123_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_16, data_out=>output_MAC_123_16);

	MAC_123_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_17, data_out=>output_MAC_123_17);

	MAC_123_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_18, data_out=>output_MAC_123_18);

	MAC_123_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_19, data_out=>output_MAC_123_19);

	MAC_123_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_20, data_out=>output_MAC_123_20);

	MAC_123_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_21, data_out=>output_MAC_123_21);

	MAC_123_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_22, data_out=>output_MAC_123_22);

	MAC_123_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_23, data_out=>output_MAC_123_23);

	MAC_123_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_24, data_out=>output_MAC_123_24);

	MAC_123_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_25, data_out=>output_MAC_123_25);

	MAC_123_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_26, data_out=>output_MAC_123_26);

	MAC_123_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_27, data_out=>output_MAC_123_27);

	MAC_123_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_28, data_out=>output_MAC_123_28);

	MAC_123_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_29, data_out=>output_MAC_123_29);

	MAC_123_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_30, data_out=>output_MAC_123_30);

	MAC_123_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_123, data_in_B=>reg_input_col_31, data_out=>output_MAC_123_31);

	MAC_124_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_0, data_out=>output_MAC_124_0);

	MAC_124_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_1, data_out=>output_MAC_124_1);

	MAC_124_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_2, data_out=>output_MAC_124_2);

	MAC_124_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_3, data_out=>output_MAC_124_3);

	MAC_124_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_4, data_out=>output_MAC_124_4);

	MAC_124_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_5, data_out=>output_MAC_124_5);

	MAC_124_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_6, data_out=>output_MAC_124_6);

	MAC_124_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_7, data_out=>output_MAC_124_7);

	MAC_124_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_8, data_out=>output_MAC_124_8);

	MAC_124_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_9, data_out=>output_MAC_124_9);

	MAC_124_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_10, data_out=>output_MAC_124_10);

	MAC_124_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_11, data_out=>output_MAC_124_11);

	MAC_124_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_12, data_out=>output_MAC_124_12);

	MAC_124_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_13, data_out=>output_MAC_124_13);

	MAC_124_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_14, data_out=>output_MAC_124_14);

	MAC_124_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_15, data_out=>output_MAC_124_15);

	MAC_124_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_16, data_out=>output_MAC_124_16);

	MAC_124_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_17, data_out=>output_MAC_124_17);

	MAC_124_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_18, data_out=>output_MAC_124_18);

	MAC_124_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_19, data_out=>output_MAC_124_19);

	MAC_124_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_20, data_out=>output_MAC_124_20);

	MAC_124_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_21, data_out=>output_MAC_124_21);

	MAC_124_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_22, data_out=>output_MAC_124_22);

	MAC_124_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_23, data_out=>output_MAC_124_23);

	MAC_124_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_24, data_out=>output_MAC_124_24);

	MAC_124_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_25, data_out=>output_MAC_124_25);

	MAC_124_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_26, data_out=>output_MAC_124_26);

	MAC_124_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_27, data_out=>output_MAC_124_27);

	MAC_124_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_28, data_out=>output_MAC_124_28);

	MAC_124_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_29, data_out=>output_MAC_124_29);

	MAC_124_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_30, data_out=>output_MAC_124_30);

	MAC_124_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_124, data_in_B=>reg_input_col_31, data_out=>output_MAC_124_31);

	MAC_125_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_0, data_out=>output_MAC_125_0);

	MAC_125_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_1, data_out=>output_MAC_125_1);

	MAC_125_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_2, data_out=>output_MAC_125_2);

	MAC_125_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_3, data_out=>output_MAC_125_3);

	MAC_125_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_4, data_out=>output_MAC_125_4);

	MAC_125_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_5, data_out=>output_MAC_125_5);

	MAC_125_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_6, data_out=>output_MAC_125_6);

	MAC_125_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_7, data_out=>output_MAC_125_7);

	MAC_125_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_8, data_out=>output_MAC_125_8);

	MAC_125_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_9, data_out=>output_MAC_125_9);

	MAC_125_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_10, data_out=>output_MAC_125_10);

	MAC_125_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_11, data_out=>output_MAC_125_11);

	MAC_125_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_12, data_out=>output_MAC_125_12);

	MAC_125_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_13, data_out=>output_MAC_125_13);

	MAC_125_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_14, data_out=>output_MAC_125_14);

	MAC_125_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_15, data_out=>output_MAC_125_15);

	MAC_125_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_16, data_out=>output_MAC_125_16);

	MAC_125_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_17, data_out=>output_MAC_125_17);

	MAC_125_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_18, data_out=>output_MAC_125_18);

	MAC_125_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_19, data_out=>output_MAC_125_19);

	MAC_125_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_20, data_out=>output_MAC_125_20);

	MAC_125_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_21, data_out=>output_MAC_125_21);

	MAC_125_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_22, data_out=>output_MAC_125_22);

	MAC_125_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_23, data_out=>output_MAC_125_23);

	MAC_125_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_24, data_out=>output_MAC_125_24);

	MAC_125_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_25, data_out=>output_MAC_125_25);

	MAC_125_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_26, data_out=>output_MAC_125_26);

	MAC_125_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_27, data_out=>output_MAC_125_27);

	MAC_125_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_28, data_out=>output_MAC_125_28);

	MAC_125_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_29, data_out=>output_MAC_125_29);

	MAC_125_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_30, data_out=>output_MAC_125_30);

	MAC_125_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_125, data_in_B=>reg_input_col_31, data_out=>output_MAC_125_31);

	MAC_126_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_0, data_out=>output_MAC_126_0);

	MAC_126_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_1, data_out=>output_MAC_126_1);

	MAC_126_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_2, data_out=>output_MAC_126_2);

	MAC_126_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_3, data_out=>output_MAC_126_3);

	MAC_126_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_4, data_out=>output_MAC_126_4);

	MAC_126_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_5, data_out=>output_MAC_126_5);

	MAC_126_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_6, data_out=>output_MAC_126_6);

	MAC_126_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_7, data_out=>output_MAC_126_7);

	MAC_126_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_8, data_out=>output_MAC_126_8);

	MAC_126_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_9, data_out=>output_MAC_126_9);

	MAC_126_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_10, data_out=>output_MAC_126_10);

	MAC_126_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_11, data_out=>output_MAC_126_11);

	MAC_126_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_12, data_out=>output_MAC_126_12);

	MAC_126_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_13, data_out=>output_MAC_126_13);

	MAC_126_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_14, data_out=>output_MAC_126_14);

	MAC_126_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_15, data_out=>output_MAC_126_15);

	MAC_126_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_16, data_out=>output_MAC_126_16);

	MAC_126_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_17, data_out=>output_MAC_126_17);

	MAC_126_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_18, data_out=>output_MAC_126_18);

	MAC_126_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_19, data_out=>output_MAC_126_19);

	MAC_126_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_20, data_out=>output_MAC_126_20);

	MAC_126_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_21, data_out=>output_MAC_126_21);

	MAC_126_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_22, data_out=>output_MAC_126_22);

	MAC_126_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_23, data_out=>output_MAC_126_23);

	MAC_126_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_24, data_out=>output_MAC_126_24);

	MAC_126_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_25, data_out=>output_MAC_126_25);

	MAC_126_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_26, data_out=>output_MAC_126_26);

	MAC_126_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_27, data_out=>output_MAC_126_27);

	MAC_126_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_28, data_out=>output_MAC_126_28);

	MAC_126_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_29, data_out=>output_MAC_126_29);

	MAC_126_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_30, data_out=>output_MAC_126_30);

	MAC_126_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_126, data_in_B=>reg_input_col_31, data_out=>output_MAC_126_31);

	MAC_127_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_0, data_out=>output_MAC_127_0);

	MAC_127_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_1, data_out=>output_MAC_127_1);

	MAC_127_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_2, data_out=>output_MAC_127_2);

	MAC_127_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_3, data_out=>output_MAC_127_3);

	MAC_127_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_4, data_out=>output_MAC_127_4);

	MAC_127_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_5, data_out=>output_MAC_127_5);

	MAC_127_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_6, data_out=>output_MAC_127_6);

	MAC_127_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_7, data_out=>output_MAC_127_7);

	MAC_127_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_8, data_out=>output_MAC_127_8);

	MAC_127_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_9, data_out=>output_MAC_127_9);

	MAC_127_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_10, data_out=>output_MAC_127_10);

	MAC_127_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_11, data_out=>output_MAC_127_11);

	MAC_127_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_12, data_out=>output_MAC_127_12);

	MAC_127_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_13, data_out=>output_MAC_127_13);

	MAC_127_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_14, data_out=>output_MAC_127_14);

	MAC_127_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_15, data_out=>output_MAC_127_15);

	MAC_127_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_16, data_out=>output_MAC_127_16);

	MAC_127_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_17, data_out=>output_MAC_127_17);

	MAC_127_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_18, data_out=>output_MAC_127_18);

	MAC_127_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_19, data_out=>output_MAC_127_19);

	MAC_127_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_20, data_out=>output_MAC_127_20);

	MAC_127_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_21, data_out=>output_MAC_127_21);

	MAC_127_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_22, data_out=>output_MAC_127_22);

	MAC_127_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_23, data_out=>output_MAC_127_23);

	MAC_127_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_24, data_out=>output_MAC_127_24);

	MAC_127_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_25, data_out=>output_MAC_127_25);

	MAC_127_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_26, data_out=>output_MAC_127_26);

	MAC_127_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_27, data_out=>output_MAC_127_27);

	MAC_127_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_28, data_out=>output_MAC_127_28);

	MAC_127_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_29, data_out=>output_MAC_127_29);

	MAC_127_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_30, data_out=>output_MAC_127_30);

	MAC_127_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_127, data_in_B=>reg_input_col_31, data_out=>output_MAC_127_31);


	mux_row_0: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_0_0, I1=>output_MAC_0_1, I2=>output_MAC_0_2, I3=>output_MAC_0_3, I4=>output_MAC_0_4, I5=>output_MAC_0_5, I6=>output_MAC_0_6, I7=>output_MAC_0_7, I8=>output_MAC_0_8, I9=>output_MAC_0_9, I10=>output_MAC_0_10, I11=>output_MAC_0_11, I12=>output_MAC_0_12, I13=>output_MAC_0_13, I14=>output_MAC_0_14, I15=>output_MAC_0_15, I16=>output_MAC_0_16, I17=>output_MAC_0_17, I18=>output_MAC_0_18, I19=>output_MAC_0_19, I20=>output_MAC_0_20, I21=>output_MAC_0_21, I22=>output_MAC_0_22, I23=>output_MAC_0_23, I24=>output_MAC_0_24, I25=>output_MAC_0_25, I26=>output_MAC_0_26, I27=>output_MAC_0_27, I28=>output_MAC_0_28, I29=>output_MAC_0_29, I30=>output_MAC_0_30, I31=>output_MAC_0_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_0);

	mux_row_1: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_1_0, I1=>output_MAC_1_1, I2=>output_MAC_1_2, I3=>output_MAC_1_3, I4=>output_MAC_1_4, I5=>output_MAC_1_5, I6=>output_MAC_1_6, I7=>output_MAC_1_7, I8=>output_MAC_1_8, I9=>output_MAC_1_9, I10=>output_MAC_1_10, I11=>output_MAC_1_11, I12=>output_MAC_1_12, I13=>output_MAC_1_13, I14=>output_MAC_1_14, I15=>output_MAC_1_15, I16=>output_MAC_1_16, I17=>output_MAC_1_17, I18=>output_MAC_1_18, I19=>output_MAC_1_19, I20=>output_MAC_1_20, I21=>output_MAC_1_21, I22=>output_MAC_1_22, I23=>output_MAC_1_23, I24=>output_MAC_1_24, I25=>output_MAC_1_25, I26=>output_MAC_1_26, I27=>output_MAC_1_27, I28=>output_MAC_1_28, I29=>output_MAC_1_29, I30=>output_MAC_1_30, I31=>output_MAC_1_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_1);

	mux_row_2: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_2_0, I1=>output_MAC_2_1, I2=>output_MAC_2_2, I3=>output_MAC_2_3, I4=>output_MAC_2_4, I5=>output_MAC_2_5, I6=>output_MAC_2_6, I7=>output_MAC_2_7, I8=>output_MAC_2_8, I9=>output_MAC_2_9, I10=>output_MAC_2_10, I11=>output_MAC_2_11, I12=>output_MAC_2_12, I13=>output_MAC_2_13, I14=>output_MAC_2_14, I15=>output_MAC_2_15, I16=>output_MAC_2_16, I17=>output_MAC_2_17, I18=>output_MAC_2_18, I19=>output_MAC_2_19, I20=>output_MAC_2_20, I21=>output_MAC_2_21, I22=>output_MAC_2_22, I23=>output_MAC_2_23, I24=>output_MAC_2_24, I25=>output_MAC_2_25, I26=>output_MAC_2_26, I27=>output_MAC_2_27, I28=>output_MAC_2_28, I29=>output_MAC_2_29, I30=>output_MAC_2_30, I31=>output_MAC_2_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_2);

	mux_row_3: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_3_0, I1=>output_MAC_3_1, I2=>output_MAC_3_2, I3=>output_MAC_3_3, I4=>output_MAC_3_4, I5=>output_MAC_3_5, I6=>output_MAC_3_6, I7=>output_MAC_3_7, I8=>output_MAC_3_8, I9=>output_MAC_3_9, I10=>output_MAC_3_10, I11=>output_MAC_3_11, I12=>output_MAC_3_12, I13=>output_MAC_3_13, I14=>output_MAC_3_14, I15=>output_MAC_3_15, I16=>output_MAC_3_16, I17=>output_MAC_3_17, I18=>output_MAC_3_18, I19=>output_MAC_3_19, I20=>output_MAC_3_20, I21=>output_MAC_3_21, I22=>output_MAC_3_22, I23=>output_MAC_3_23, I24=>output_MAC_3_24, I25=>output_MAC_3_25, I26=>output_MAC_3_26, I27=>output_MAC_3_27, I28=>output_MAC_3_28, I29=>output_MAC_3_29, I30=>output_MAC_3_30, I31=>output_MAC_3_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_3);

	mux_row_4: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_4_0, I1=>output_MAC_4_1, I2=>output_MAC_4_2, I3=>output_MAC_4_3, I4=>output_MAC_4_4, I5=>output_MAC_4_5, I6=>output_MAC_4_6, I7=>output_MAC_4_7, I8=>output_MAC_4_8, I9=>output_MAC_4_9, I10=>output_MAC_4_10, I11=>output_MAC_4_11, I12=>output_MAC_4_12, I13=>output_MAC_4_13, I14=>output_MAC_4_14, I15=>output_MAC_4_15, I16=>output_MAC_4_16, I17=>output_MAC_4_17, I18=>output_MAC_4_18, I19=>output_MAC_4_19, I20=>output_MAC_4_20, I21=>output_MAC_4_21, I22=>output_MAC_4_22, I23=>output_MAC_4_23, I24=>output_MAC_4_24, I25=>output_MAC_4_25, I26=>output_MAC_4_26, I27=>output_MAC_4_27, I28=>output_MAC_4_28, I29=>output_MAC_4_29, I30=>output_MAC_4_30, I31=>output_MAC_4_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_4);

	mux_row_5: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_5_0, I1=>output_MAC_5_1, I2=>output_MAC_5_2, I3=>output_MAC_5_3, I4=>output_MAC_5_4, I5=>output_MAC_5_5, I6=>output_MAC_5_6, I7=>output_MAC_5_7, I8=>output_MAC_5_8, I9=>output_MAC_5_9, I10=>output_MAC_5_10, I11=>output_MAC_5_11, I12=>output_MAC_5_12, I13=>output_MAC_5_13, I14=>output_MAC_5_14, I15=>output_MAC_5_15, I16=>output_MAC_5_16, I17=>output_MAC_5_17, I18=>output_MAC_5_18, I19=>output_MAC_5_19, I20=>output_MAC_5_20, I21=>output_MAC_5_21, I22=>output_MAC_5_22, I23=>output_MAC_5_23, I24=>output_MAC_5_24, I25=>output_MAC_5_25, I26=>output_MAC_5_26, I27=>output_MAC_5_27, I28=>output_MAC_5_28, I29=>output_MAC_5_29, I30=>output_MAC_5_30, I31=>output_MAC_5_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_5);

	mux_row_6: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_6_0, I1=>output_MAC_6_1, I2=>output_MAC_6_2, I3=>output_MAC_6_3, I4=>output_MAC_6_4, I5=>output_MAC_6_5, I6=>output_MAC_6_6, I7=>output_MAC_6_7, I8=>output_MAC_6_8, I9=>output_MAC_6_9, I10=>output_MAC_6_10, I11=>output_MAC_6_11, I12=>output_MAC_6_12, I13=>output_MAC_6_13, I14=>output_MAC_6_14, I15=>output_MAC_6_15, I16=>output_MAC_6_16, I17=>output_MAC_6_17, I18=>output_MAC_6_18, I19=>output_MAC_6_19, I20=>output_MAC_6_20, I21=>output_MAC_6_21, I22=>output_MAC_6_22, I23=>output_MAC_6_23, I24=>output_MAC_6_24, I25=>output_MAC_6_25, I26=>output_MAC_6_26, I27=>output_MAC_6_27, I28=>output_MAC_6_28, I29=>output_MAC_6_29, I30=>output_MAC_6_30, I31=>output_MAC_6_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_6);

	mux_row_7: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_7_0, I1=>output_MAC_7_1, I2=>output_MAC_7_2, I3=>output_MAC_7_3, I4=>output_MAC_7_4, I5=>output_MAC_7_5, I6=>output_MAC_7_6, I7=>output_MAC_7_7, I8=>output_MAC_7_8, I9=>output_MAC_7_9, I10=>output_MAC_7_10, I11=>output_MAC_7_11, I12=>output_MAC_7_12, I13=>output_MAC_7_13, I14=>output_MAC_7_14, I15=>output_MAC_7_15, I16=>output_MAC_7_16, I17=>output_MAC_7_17, I18=>output_MAC_7_18, I19=>output_MAC_7_19, I20=>output_MAC_7_20, I21=>output_MAC_7_21, I22=>output_MAC_7_22, I23=>output_MAC_7_23, I24=>output_MAC_7_24, I25=>output_MAC_7_25, I26=>output_MAC_7_26, I27=>output_MAC_7_27, I28=>output_MAC_7_28, I29=>output_MAC_7_29, I30=>output_MAC_7_30, I31=>output_MAC_7_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_7);

	mux_row_8: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_8_0, I1=>output_MAC_8_1, I2=>output_MAC_8_2, I3=>output_MAC_8_3, I4=>output_MAC_8_4, I5=>output_MAC_8_5, I6=>output_MAC_8_6, I7=>output_MAC_8_7, I8=>output_MAC_8_8, I9=>output_MAC_8_9, I10=>output_MAC_8_10, I11=>output_MAC_8_11, I12=>output_MAC_8_12, I13=>output_MAC_8_13, I14=>output_MAC_8_14, I15=>output_MAC_8_15, I16=>output_MAC_8_16, I17=>output_MAC_8_17, I18=>output_MAC_8_18, I19=>output_MAC_8_19, I20=>output_MAC_8_20, I21=>output_MAC_8_21, I22=>output_MAC_8_22, I23=>output_MAC_8_23, I24=>output_MAC_8_24, I25=>output_MAC_8_25, I26=>output_MAC_8_26, I27=>output_MAC_8_27, I28=>output_MAC_8_28, I29=>output_MAC_8_29, I30=>output_MAC_8_30, I31=>output_MAC_8_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_8);

	mux_row_9: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_9_0, I1=>output_MAC_9_1, I2=>output_MAC_9_2, I3=>output_MAC_9_3, I4=>output_MAC_9_4, I5=>output_MAC_9_5, I6=>output_MAC_9_6, I7=>output_MAC_9_7, I8=>output_MAC_9_8, I9=>output_MAC_9_9, I10=>output_MAC_9_10, I11=>output_MAC_9_11, I12=>output_MAC_9_12, I13=>output_MAC_9_13, I14=>output_MAC_9_14, I15=>output_MAC_9_15, I16=>output_MAC_9_16, I17=>output_MAC_9_17, I18=>output_MAC_9_18, I19=>output_MAC_9_19, I20=>output_MAC_9_20, I21=>output_MAC_9_21, I22=>output_MAC_9_22, I23=>output_MAC_9_23, I24=>output_MAC_9_24, I25=>output_MAC_9_25, I26=>output_MAC_9_26, I27=>output_MAC_9_27, I28=>output_MAC_9_28, I29=>output_MAC_9_29, I30=>output_MAC_9_30, I31=>output_MAC_9_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_9);

	mux_row_10: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_10_0, I1=>output_MAC_10_1, I2=>output_MAC_10_2, I3=>output_MAC_10_3, I4=>output_MAC_10_4, I5=>output_MAC_10_5, I6=>output_MAC_10_6, I7=>output_MAC_10_7, I8=>output_MAC_10_8, I9=>output_MAC_10_9, I10=>output_MAC_10_10, I11=>output_MAC_10_11, I12=>output_MAC_10_12, I13=>output_MAC_10_13, I14=>output_MAC_10_14, I15=>output_MAC_10_15, I16=>output_MAC_10_16, I17=>output_MAC_10_17, I18=>output_MAC_10_18, I19=>output_MAC_10_19, I20=>output_MAC_10_20, I21=>output_MAC_10_21, I22=>output_MAC_10_22, I23=>output_MAC_10_23, I24=>output_MAC_10_24, I25=>output_MAC_10_25, I26=>output_MAC_10_26, I27=>output_MAC_10_27, I28=>output_MAC_10_28, I29=>output_MAC_10_29, I30=>output_MAC_10_30, I31=>output_MAC_10_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_10);

	mux_row_11: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_11_0, I1=>output_MAC_11_1, I2=>output_MAC_11_2, I3=>output_MAC_11_3, I4=>output_MAC_11_4, I5=>output_MAC_11_5, I6=>output_MAC_11_6, I7=>output_MAC_11_7, I8=>output_MAC_11_8, I9=>output_MAC_11_9, I10=>output_MAC_11_10, I11=>output_MAC_11_11, I12=>output_MAC_11_12, I13=>output_MAC_11_13, I14=>output_MAC_11_14, I15=>output_MAC_11_15, I16=>output_MAC_11_16, I17=>output_MAC_11_17, I18=>output_MAC_11_18, I19=>output_MAC_11_19, I20=>output_MAC_11_20, I21=>output_MAC_11_21, I22=>output_MAC_11_22, I23=>output_MAC_11_23, I24=>output_MAC_11_24, I25=>output_MAC_11_25, I26=>output_MAC_11_26, I27=>output_MAC_11_27, I28=>output_MAC_11_28, I29=>output_MAC_11_29, I30=>output_MAC_11_30, I31=>output_MAC_11_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_11);

	mux_row_12: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_12_0, I1=>output_MAC_12_1, I2=>output_MAC_12_2, I3=>output_MAC_12_3, I4=>output_MAC_12_4, I5=>output_MAC_12_5, I6=>output_MAC_12_6, I7=>output_MAC_12_7, I8=>output_MAC_12_8, I9=>output_MAC_12_9, I10=>output_MAC_12_10, I11=>output_MAC_12_11, I12=>output_MAC_12_12, I13=>output_MAC_12_13, I14=>output_MAC_12_14, I15=>output_MAC_12_15, I16=>output_MAC_12_16, I17=>output_MAC_12_17, I18=>output_MAC_12_18, I19=>output_MAC_12_19, I20=>output_MAC_12_20, I21=>output_MAC_12_21, I22=>output_MAC_12_22, I23=>output_MAC_12_23, I24=>output_MAC_12_24, I25=>output_MAC_12_25, I26=>output_MAC_12_26, I27=>output_MAC_12_27, I28=>output_MAC_12_28, I29=>output_MAC_12_29, I30=>output_MAC_12_30, I31=>output_MAC_12_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_12);

	mux_row_13: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_13_0, I1=>output_MAC_13_1, I2=>output_MAC_13_2, I3=>output_MAC_13_3, I4=>output_MAC_13_4, I5=>output_MAC_13_5, I6=>output_MAC_13_6, I7=>output_MAC_13_7, I8=>output_MAC_13_8, I9=>output_MAC_13_9, I10=>output_MAC_13_10, I11=>output_MAC_13_11, I12=>output_MAC_13_12, I13=>output_MAC_13_13, I14=>output_MAC_13_14, I15=>output_MAC_13_15, I16=>output_MAC_13_16, I17=>output_MAC_13_17, I18=>output_MAC_13_18, I19=>output_MAC_13_19, I20=>output_MAC_13_20, I21=>output_MAC_13_21, I22=>output_MAC_13_22, I23=>output_MAC_13_23, I24=>output_MAC_13_24, I25=>output_MAC_13_25, I26=>output_MAC_13_26, I27=>output_MAC_13_27, I28=>output_MAC_13_28, I29=>output_MAC_13_29, I30=>output_MAC_13_30, I31=>output_MAC_13_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_13);

	mux_row_14: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_14_0, I1=>output_MAC_14_1, I2=>output_MAC_14_2, I3=>output_MAC_14_3, I4=>output_MAC_14_4, I5=>output_MAC_14_5, I6=>output_MAC_14_6, I7=>output_MAC_14_7, I8=>output_MAC_14_8, I9=>output_MAC_14_9, I10=>output_MAC_14_10, I11=>output_MAC_14_11, I12=>output_MAC_14_12, I13=>output_MAC_14_13, I14=>output_MAC_14_14, I15=>output_MAC_14_15, I16=>output_MAC_14_16, I17=>output_MAC_14_17, I18=>output_MAC_14_18, I19=>output_MAC_14_19, I20=>output_MAC_14_20, I21=>output_MAC_14_21, I22=>output_MAC_14_22, I23=>output_MAC_14_23, I24=>output_MAC_14_24, I25=>output_MAC_14_25, I26=>output_MAC_14_26, I27=>output_MAC_14_27, I28=>output_MAC_14_28, I29=>output_MAC_14_29, I30=>output_MAC_14_30, I31=>output_MAC_14_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_14);

	mux_row_15: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_15_0, I1=>output_MAC_15_1, I2=>output_MAC_15_2, I3=>output_MAC_15_3, I4=>output_MAC_15_4, I5=>output_MAC_15_5, I6=>output_MAC_15_6, I7=>output_MAC_15_7, I8=>output_MAC_15_8, I9=>output_MAC_15_9, I10=>output_MAC_15_10, I11=>output_MAC_15_11, I12=>output_MAC_15_12, I13=>output_MAC_15_13, I14=>output_MAC_15_14, I15=>output_MAC_15_15, I16=>output_MAC_15_16, I17=>output_MAC_15_17, I18=>output_MAC_15_18, I19=>output_MAC_15_19, I20=>output_MAC_15_20, I21=>output_MAC_15_21, I22=>output_MAC_15_22, I23=>output_MAC_15_23, I24=>output_MAC_15_24, I25=>output_MAC_15_25, I26=>output_MAC_15_26, I27=>output_MAC_15_27, I28=>output_MAC_15_28, I29=>output_MAC_15_29, I30=>output_MAC_15_30, I31=>output_MAC_15_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_15);

	mux_row_16: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_16_0, I1=>output_MAC_16_1, I2=>output_MAC_16_2, I3=>output_MAC_16_3, I4=>output_MAC_16_4, I5=>output_MAC_16_5, I6=>output_MAC_16_6, I7=>output_MAC_16_7, I8=>output_MAC_16_8, I9=>output_MAC_16_9, I10=>output_MAC_16_10, I11=>output_MAC_16_11, I12=>output_MAC_16_12, I13=>output_MAC_16_13, I14=>output_MAC_16_14, I15=>output_MAC_16_15, I16=>output_MAC_16_16, I17=>output_MAC_16_17, I18=>output_MAC_16_18, I19=>output_MAC_16_19, I20=>output_MAC_16_20, I21=>output_MAC_16_21, I22=>output_MAC_16_22, I23=>output_MAC_16_23, I24=>output_MAC_16_24, I25=>output_MAC_16_25, I26=>output_MAC_16_26, I27=>output_MAC_16_27, I28=>output_MAC_16_28, I29=>output_MAC_16_29, I30=>output_MAC_16_30, I31=>output_MAC_16_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_16);

	mux_row_17: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_17_0, I1=>output_MAC_17_1, I2=>output_MAC_17_2, I3=>output_MAC_17_3, I4=>output_MAC_17_4, I5=>output_MAC_17_5, I6=>output_MAC_17_6, I7=>output_MAC_17_7, I8=>output_MAC_17_8, I9=>output_MAC_17_9, I10=>output_MAC_17_10, I11=>output_MAC_17_11, I12=>output_MAC_17_12, I13=>output_MAC_17_13, I14=>output_MAC_17_14, I15=>output_MAC_17_15, I16=>output_MAC_17_16, I17=>output_MAC_17_17, I18=>output_MAC_17_18, I19=>output_MAC_17_19, I20=>output_MAC_17_20, I21=>output_MAC_17_21, I22=>output_MAC_17_22, I23=>output_MAC_17_23, I24=>output_MAC_17_24, I25=>output_MAC_17_25, I26=>output_MAC_17_26, I27=>output_MAC_17_27, I28=>output_MAC_17_28, I29=>output_MAC_17_29, I30=>output_MAC_17_30, I31=>output_MAC_17_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_17);

	mux_row_18: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_18_0, I1=>output_MAC_18_1, I2=>output_MAC_18_2, I3=>output_MAC_18_3, I4=>output_MAC_18_4, I5=>output_MAC_18_5, I6=>output_MAC_18_6, I7=>output_MAC_18_7, I8=>output_MAC_18_8, I9=>output_MAC_18_9, I10=>output_MAC_18_10, I11=>output_MAC_18_11, I12=>output_MAC_18_12, I13=>output_MAC_18_13, I14=>output_MAC_18_14, I15=>output_MAC_18_15, I16=>output_MAC_18_16, I17=>output_MAC_18_17, I18=>output_MAC_18_18, I19=>output_MAC_18_19, I20=>output_MAC_18_20, I21=>output_MAC_18_21, I22=>output_MAC_18_22, I23=>output_MAC_18_23, I24=>output_MAC_18_24, I25=>output_MAC_18_25, I26=>output_MAC_18_26, I27=>output_MAC_18_27, I28=>output_MAC_18_28, I29=>output_MAC_18_29, I30=>output_MAC_18_30, I31=>output_MAC_18_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_18);

	mux_row_19: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_19_0, I1=>output_MAC_19_1, I2=>output_MAC_19_2, I3=>output_MAC_19_3, I4=>output_MAC_19_4, I5=>output_MAC_19_5, I6=>output_MAC_19_6, I7=>output_MAC_19_7, I8=>output_MAC_19_8, I9=>output_MAC_19_9, I10=>output_MAC_19_10, I11=>output_MAC_19_11, I12=>output_MAC_19_12, I13=>output_MAC_19_13, I14=>output_MAC_19_14, I15=>output_MAC_19_15, I16=>output_MAC_19_16, I17=>output_MAC_19_17, I18=>output_MAC_19_18, I19=>output_MAC_19_19, I20=>output_MAC_19_20, I21=>output_MAC_19_21, I22=>output_MAC_19_22, I23=>output_MAC_19_23, I24=>output_MAC_19_24, I25=>output_MAC_19_25, I26=>output_MAC_19_26, I27=>output_MAC_19_27, I28=>output_MAC_19_28, I29=>output_MAC_19_29, I30=>output_MAC_19_30, I31=>output_MAC_19_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_19);

	mux_row_20: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_20_0, I1=>output_MAC_20_1, I2=>output_MAC_20_2, I3=>output_MAC_20_3, I4=>output_MAC_20_4, I5=>output_MAC_20_5, I6=>output_MAC_20_6, I7=>output_MAC_20_7, I8=>output_MAC_20_8, I9=>output_MAC_20_9, I10=>output_MAC_20_10, I11=>output_MAC_20_11, I12=>output_MAC_20_12, I13=>output_MAC_20_13, I14=>output_MAC_20_14, I15=>output_MAC_20_15, I16=>output_MAC_20_16, I17=>output_MAC_20_17, I18=>output_MAC_20_18, I19=>output_MAC_20_19, I20=>output_MAC_20_20, I21=>output_MAC_20_21, I22=>output_MAC_20_22, I23=>output_MAC_20_23, I24=>output_MAC_20_24, I25=>output_MAC_20_25, I26=>output_MAC_20_26, I27=>output_MAC_20_27, I28=>output_MAC_20_28, I29=>output_MAC_20_29, I30=>output_MAC_20_30, I31=>output_MAC_20_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_20);

	mux_row_21: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_21_0, I1=>output_MAC_21_1, I2=>output_MAC_21_2, I3=>output_MAC_21_3, I4=>output_MAC_21_4, I5=>output_MAC_21_5, I6=>output_MAC_21_6, I7=>output_MAC_21_7, I8=>output_MAC_21_8, I9=>output_MAC_21_9, I10=>output_MAC_21_10, I11=>output_MAC_21_11, I12=>output_MAC_21_12, I13=>output_MAC_21_13, I14=>output_MAC_21_14, I15=>output_MAC_21_15, I16=>output_MAC_21_16, I17=>output_MAC_21_17, I18=>output_MAC_21_18, I19=>output_MAC_21_19, I20=>output_MAC_21_20, I21=>output_MAC_21_21, I22=>output_MAC_21_22, I23=>output_MAC_21_23, I24=>output_MAC_21_24, I25=>output_MAC_21_25, I26=>output_MAC_21_26, I27=>output_MAC_21_27, I28=>output_MAC_21_28, I29=>output_MAC_21_29, I30=>output_MAC_21_30, I31=>output_MAC_21_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_21);

	mux_row_22: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_22_0, I1=>output_MAC_22_1, I2=>output_MAC_22_2, I3=>output_MAC_22_3, I4=>output_MAC_22_4, I5=>output_MAC_22_5, I6=>output_MAC_22_6, I7=>output_MAC_22_7, I8=>output_MAC_22_8, I9=>output_MAC_22_9, I10=>output_MAC_22_10, I11=>output_MAC_22_11, I12=>output_MAC_22_12, I13=>output_MAC_22_13, I14=>output_MAC_22_14, I15=>output_MAC_22_15, I16=>output_MAC_22_16, I17=>output_MAC_22_17, I18=>output_MAC_22_18, I19=>output_MAC_22_19, I20=>output_MAC_22_20, I21=>output_MAC_22_21, I22=>output_MAC_22_22, I23=>output_MAC_22_23, I24=>output_MAC_22_24, I25=>output_MAC_22_25, I26=>output_MAC_22_26, I27=>output_MAC_22_27, I28=>output_MAC_22_28, I29=>output_MAC_22_29, I30=>output_MAC_22_30, I31=>output_MAC_22_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_22);

	mux_row_23: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_23_0, I1=>output_MAC_23_1, I2=>output_MAC_23_2, I3=>output_MAC_23_3, I4=>output_MAC_23_4, I5=>output_MAC_23_5, I6=>output_MAC_23_6, I7=>output_MAC_23_7, I8=>output_MAC_23_8, I9=>output_MAC_23_9, I10=>output_MAC_23_10, I11=>output_MAC_23_11, I12=>output_MAC_23_12, I13=>output_MAC_23_13, I14=>output_MAC_23_14, I15=>output_MAC_23_15, I16=>output_MAC_23_16, I17=>output_MAC_23_17, I18=>output_MAC_23_18, I19=>output_MAC_23_19, I20=>output_MAC_23_20, I21=>output_MAC_23_21, I22=>output_MAC_23_22, I23=>output_MAC_23_23, I24=>output_MAC_23_24, I25=>output_MAC_23_25, I26=>output_MAC_23_26, I27=>output_MAC_23_27, I28=>output_MAC_23_28, I29=>output_MAC_23_29, I30=>output_MAC_23_30, I31=>output_MAC_23_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_23);

	mux_row_24: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_24_0, I1=>output_MAC_24_1, I2=>output_MAC_24_2, I3=>output_MAC_24_3, I4=>output_MAC_24_4, I5=>output_MAC_24_5, I6=>output_MAC_24_6, I7=>output_MAC_24_7, I8=>output_MAC_24_8, I9=>output_MAC_24_9, I10=>output_MAC_24_10, I11=>output_MAC_24_11, I12=>output_MAC_24_12, I13=>output_MAC_24_13, I14=>output_MAC_24_14, I15=>output_MAC_24_15, I16=>output_MAC_24_16, I17=>output_MAC_24_17, I18=>output_MAC_24_18, I19=>output_MAC_24_19, I20=>output_MAC_24_20, I21=>output_MAC_24_21, I22=>output_MAC_24_22, I23=>output_MAC_24_23, I24=>output_MAC_24_24, I25=>output_MAC_24_25, I26=>output_MAC_24_26, I27=>output_MAC_24_27, I28=>output_MAC_24_28, I29=>output_MAC_24_29, I30=>output_MAC_24_30, I31=>output_MAC_24_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_24);

	mux_row_25: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_25_0, I1=>output_MAC_25_1, I2=>output_MAC_25_2, I3=>output_MAC_25_3, I4=>output_MAC_25_4, I5=>output_MAC_25_5, I6=>output_MAC_25_6, I7=>output_MAC_25_7, I8=>output_MAC_25_8, I9=>output_MAC_25_9, I10=>output_MAC_25_10, I11=>output_MAC_25_11, I12=>output_MAC_25_12, I13=>output_MAC_25_13, I14=>output_MAC_25_14, I15=>output_MAC_25_15, I16=>output_MAC_25_16, I17=>output_MAC_25_17, I18=>output_MAC_25_18, I19=>output_MAC_25_19, I20=>output_MAC_25_20, I21=>output_MAC_25_21, I22=>output_MAC_25_22, I23=>output_MAC_25_23, I24=>output_MAC_25_24, I25=>output_MAC_25_25, I26=>output_MAC_25_26, I27=>output_MAC_25_27, I28=>output_MAC_25_28, I29=>output_MAC_25_29, I30=>output_MAC_25_30, I31=>output_MAC_25_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_25);

	mux_row_26: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_26_0, I1=>output_MAC_26_1, I2=>output_MAC_26_2, I3=>output_MAC_26_3, I4=>output_MAC_26_4, I5=>output_MAC_26_5, I6=>output_MAC_26_6, I7=>output_MAC_26_7, I8=>output_MAC_26_8, I9=>output_MAC_26_9, I10=>output_MAC_26_10, I11=>output_MAC_26_11, I12=>output_MAC_26_12, I13=>output_MAC_26_13, I14=>output_MAC_26_14, I15=>output_MAC_26_15, I16=>output_MAC_26_16, I17=>output_MAC_26_17, I18=>output_MAC_26_18, I19=>output_MAC_26_19, I20=>output_MAC_26_20, I21=>output_MAC_26_21, I22=>output_MAC_26_22, I23=>output_MAC_26_23, I24=>output_MAC_26_24, I25=>output_MAC_26_25, I26=>output_MAC_26_26, I27=>output_MAC_26_27, I28=>output_MAC_26_28, I29=>output_MAC_26_29, I30=>output_MAC_26_30, I31=>output_MAC_26_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_26);

	mux_row_27: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_27_0, I1=>output_MAC_27_1, I2=>output_MAC_27_2, I3=>output_MAC_27_3, I4=>output_MAC_27_4, I5=>output_MAC_27_5, I6=>output_MAC_27_6, I7=>output_MAC_27_7, I8=>output_MAC_27_8, I9=>output_MAC_27_9, I10=>output_MAC_27_10, I11=>output_MAC_27_11, I12=>output_MAC_27_12, I13=>output_MAC_27_13, I14=>output_MAC_27_14, I15=>output_MAC_27_15, I16=>output_MAC_27_16, I17=>output_MAC_27_17, I18=>output_MAC_27_18, I19=>output_MAC_27_19, I20=>output_MAC_27_20, I21=>output_MAC_27_21, I22=>output_MAC_27_22, I23=>output_MAC_27_23, I24=>output_MAC_27_24, I25=>output_MAC_27_25, I26=>output_MAC_27_26, I27=>output_MAC_27_27, I28=>output_MAC_27_28, I29=>output_MAC_27_29, I30=>output_MAC_27_30, I31=>output_MAC_27_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_27);

	mux_row_28: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_28_0, I1=>output_MAC_28_1, I2=>output_MAC_28_2, I3=>output_MAC_28_3, I4=>output_MAC_28_4, I5=>output_MAC_28_5, I6=>output_MAC_28_6, I7=>output_MAC_28_7, I8=>output_MAC_28_8, I9=>output_MAC_28_9, I10=>output_MAC_28_10, I11=>output_MAC_28_11, I12=>output_MAC_28_12, I13=>output_MAC_28_13, I14=>output_MAC_28_14, I15=>output_MAC_28_15, I16=>output_MAC_28_16, I17=>output_MAC_28_17, I18=>output_MAC_28_18, I19=>output_MAC_28_19, I20=>output_MAC_28_20, I21=>output_MAC_28_21, I22=>output_MAC_28_22, I23=>output_MAC_28_23, I24=>output_MAC_28_24, I25=>output_MAC_28_25, I26=>output_MAC_28_26, I27=>output_MAC_28_27, I28=>output_MAC_28_28, I29=>output_MAC_28_29, I30=>output_MAC_28_30, I31=>output_MAC_28_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_28);

	mux_row_29: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_29_0, I1=>output_MAC_29_1, I2=>output_MAC_29_2, I3=>output_MAC_29_3, I4=>output_MAC_29_4, I5=>output_MAC_29_5, I6=>output_MAC_29_6, I7=>output_MAC_29_7, I8=>output_MAC_29_8, I9=>output_MAC_29_9, I10=>output_MAC_29_10, I11=>output_MAC_29_11, I12=>output_MAC_29_12, I13=>output_MAC_29_13, I14=>output_MAC_29_14, I15=>output_MAC_29_15, I16=>output_MAC_29_16, I17=>output_MAC_29_17, I18=>output_MAC_29_18, I19=>output_MAC_29_19, I20=>output_MAC_29_20, I21=>output_MAC_29_21, I22=>output_MAC_29_22, I23=>output_MAC_29_23, I24=>output_MAC_29_24, I25=>output_MAC_29_25, I26=>output_MAC_29_26, I27=>output_MAC_29_27, I28=>output_MAC_29_28, I29=>output_MAC_29_29, I30=>output_MAC_29_30, I31=>output_MAC_29_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_29);

	mux_row_30: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_30_0, I1=>output_MAC_30_1, I2=>output_MAC_30_2, I3=>output_MAC_30_3, I4=>output_MAC_30_4, I5=>output_MAC_30_5, I6=>output_MAC_30_6, I7=>output_MAC_30_7, I8=>output_MAC_30_8, I9=>output_MAC_30_9, I10=>output_MAC_30_10, I11=>output_MAC_30_11, I12=>output_MAC_30_12, I13=>output_MAC_30_13, I14=>output_MAC_30_14, I15=>output_MAC_30_15, I16=>output_MAC_30_16, I17=>output_MAC_30_17, I18=>output_MAC_30_18, I19=>output_MAC_30_19, I20=>output_MAC_30_20, I21=>output_MAC_30_21, I22=>output_MAC_30_22, I23=>output_MAC_30_23, I24=>output_MAC_30_24, I25=>output_MAC_30_25, I26=>output_MAC_30_26, I27=>output_MAC_30_27, I28=>output_MAC_30_28, I29=>output_MAC_30_29, I30=>output_MAC_30_30, I31=>output_MAC_30_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_30);

	mux_row_31: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_31_0, I1=>output_MAC_31_1, I2=>output_MAC_31_2, I3=>output_MAC_31_3, I4=>output_MAC_31_4, I5=>output_MAC_31_5, I6=>output_MAC_31_6, I7=>output_MAC_31_7, I8=>output_MAC_31_8, I9=>output_MAC_31_9, I10=>output_MAC_31_10, I11=>output_MAC_31_11, I12=>output_MAC_31_12, I13=>output_MAC_31_13, I14=>output_MAC_31_14, I15=>output_MAC_31_15, I16=>output_MAC_31_16, I17=>output_MAC_31_17, I18=>output_MAC_31_18, I19=>output_MAC_31_19, I20=>output_MAC_31_20, I21=>output_MAC_31_21, I22=>output_MAC_31_22, I23=>output_MAC_31_23, I24=>output_MAC_31_24, I25=>output_MAC_31_25, I26=>output_MAC_31_26, I27=>output_MAC_31_27, I28=>output_MAC_31_28, I29=>output_MAC_31_29, I30=>output_MAC_31_30, I31=>output_MAC_31_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_31);

	mux_row_32: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_32_0, I1=>output_MAC_32_1, I2=>output_MAC_32_2, I3=>output_MAC_32_3, I4=>output_MAC_32_4, I5=>output_MAC_32_5, I6=>output_MAC_32_6, I7=>output_MAC_32_7, I8=>output_MAC_32_8, I9=>output_MAC_32_9, I10=>output_MAC_32_10, I11=>output_MAC_32_11, I12=>output_MAC_32_12, I13=>output_MAC_32_13, I14=>output_MAC_32_14, I15=>output_MAC_32_15, I16=>output_MAC_32_16, I17=>output_MAC_32_17, I18=>output_MAC_32_18, I19=>output_MAC_32_19, I20=>output_MAC_32_20, I21=>output_MAC_32_21, I22=>output_MAC_32_22, I23=>output_MAC_32_23, I24=>output_MAC_32_24, I25=>output_MAC_32_25, I26=>output_MAC_32_26, I27=>output_MAC_32_27, I28=>output_MAC_32_28, I29=>output_MAC_32_29, I30=>output_MAC_32_30, I31=>output_MAC_32_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_32);

	mux_row_33: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_33_0, I1=>output_MAC_33_1, I2=>output_MAC_33_2, I3=>output_MAC_33_3, I4=>output_MAC_33_4, I5=>output_MAC_33_5, I6=>output_MAC_33_6, I7=>output_MAC_33_7, I8=>output_MAC_33_8, I9=>output_MAC_33_9, I10=>output_MAC_33_10, I11=>output_MAC_33_11, I12=>output_MAC_33_12, I13=>output_MAC_33_13, I14=>output_MAC_33_14, I15=>output_MAC_33_15, I16=>output_MAC_33_16, I17=>output_MAC_33_17, I18=>output_MAC_33_18, I19=>output_MAC_33_19, I20=>output_MAC_33_20, I21=>output_MAC_33_21, I22=>output_MAC_33_22, I23=>output_MAC_33_23, I24=>output_MAC_33_24, I25=>output_MAC_33_25, I26=>output_MAC_33_26, I27=>output_MAC_33_27, I28=>output_MAC_33_28, I29=>output_MAC_33_29, I30=>output_MAC_33_30, I31=>output_MAC_33_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_33);

	mux_row_34: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_34_0, I1=>output_MAC_34_1, I2=>output_MAC_34_2, I3=>output_MAC_34_3, I4=>output_MAC_34_4, I5=>output_MAC_34_5, I6=>output_MAC_34_6, I7=>output_MAC_34_7, I8=>output_MAC_34_8, I9=>output_MAC_34_9, I10=>output_MAC_34_10, I11=>output_MAC_34_11, I12=>output_MAC_34_12, I13=>output_MAC_34_13, I14=>output_MAC_34_14, I15=>output_MAC_34_15, I16=>output_MAC_34_16, I17=>output_MAC_34_17, I18=>output_MAC_34_18, I19=>output_MAC_34_19, I20=>output_MAC_34_20, I21=>output_MAC_34_21, I22=>output_MAC_34_22, I23=>output_MAC_34_23, I24=>output_MAC_34_24, I25=>output_MAC_34_25, I26=>output_MAC_34_26, I27=>output_MAC_34_27, I28=>output_MAC_34_28, I29=>output_MAC_34_29, I30=>output_MAC_34_30, I31=>output_MAC_34_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_34);

	mux_row_35: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_35_0, I1=>output_MAC_35_1, I2=>output_MAC_35_2, I3=>output_MAC_35_3, I4=>output_MAC_35_4, I5=>output_MAC_35_5, I6=>output_MAC_35_6, I7=>output_MAC_35_7, I8=>output_MAC_35_8, I9=>output_MAC_35_9, I10=>output_MAC_35_10, I11=>output_MAC_35_11, I12=>output_MAC_35_12, I13=>output_MAC_35_13, I14=>output_MAC_35_14, I15=>output_MAC_35_15, I16=>output_MAC_35_16, I17=>output_MAC_35_17, I18=>output_MAC_35_18, I19=>output_MAC_35_19, I20=>output_MAC_35_20, I21=>output_MAC_35_21, I22=>output_MAC_35_22, I23=>output_MAC_35_23, I24=>output_MAC_35_24, I25=>output_MAC_35_25, I26=>output_MAC_35_26, I27=>output_MAC_35_27, I28=>output_MAC_35_28, I29=>output_MAC_35_29, I30=>output_MAC_35_30, I31=>output_MAC_35_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_35);

	mux_row_36: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_36_0, I1=>output_MAC_36_1, I2=>output_MAC_36_2, I3=>output_MAC_36_3, I4=>output_MAC_36_4, I5=>output_MAC_36_5, I6=>output_MAC_36_6, I7=>output_MAC_36_7, I8=>output_MAC_36_8, I9=>output_MAC_36_9, I10=>output_MAC_36_10, I11=>output_MAC_36_11, I12=>output_MAC_36_12, I13=>output_MAC_36_13, I14=>output_MAC_36_14, I15=>output_MAC_36_15, I16=>output_MAC_36_16, I17=>output_MAC_36_17, I18=>output_MAC_36_18, I19=>output_MAC_36_19, I20=>output_MAC_36_20, I21=>output_MAC_36_21, I22=>output_MAC_36_22, I23=>output_MAC_36_23, I24=>output_MAC_36_24, I25=>output_MAC_36_25, I26=>output_MAC_36_26, I27=>output_MAC_36_27, I28=>output_MAC_36_28, I29=>output_MAC_36_29, I30=>output_MAC_36_30, I31=>output_MAC_36_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_36);

	mux_row_37: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_37_0, I1=>output_MAC_37_1, I2=>output_MAC_37_2, I3=>output_MAC_37_3, I4=>output_MAC_37_4, I5=>output_MAC_37_5, I6=>output_MAC_37_6, I7=>output_MAC_37_7, I8=>output_MAC_37_8, I9=>output_MAC_37_9, I10=>output_MAC_37_10, I11=>output_MAC_37_11, I12=>output_MAC_37_12, I13=>output_MAC_37_13, I14=>output_MAC_37_14, I15=>output_MAC_37_15, I16=>output_MAC_37_16, I17=>output_MAC_37_17, I18=>output_MAC_37_18, I19=>output_MAC_37_19, I20=>output_MAC_37_20, I21=>output_MAC_37_21, I22=>output_MAC_37_22, I23=>output_MAC_37_23, I24=>output_MAC_37_24, I25=>output_MAC_37_25, I26=>output_MAC_37_26, I27=>output_MAC_37_27, I28=>output_MAC_37_28, I29=>output_MAC_37_29, I30=>output_MAC_37_30, I31=>output_MAC_37_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_37);

	mux_row_38: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_38_0, I1=>output_MAC_38_1, I2=>output_MAC_38_2, I3=>output_MAC_38_3, I4=>output_MAC_38_4, I5=>output_MAC_38_5, I6=>output_MAC_38_6, I7=>output_MAC_38_7, I8=>output_MAC_38_8, I9=>output_MAC_38_9, I10=>output_MAC_38_10, I11=>output_MAC_38_11, I12=>output_MAC_38_12, I13=>output_MAC_38_13, I14=>output_MAC_38_14, I15=>output_MAC_38_15, I16=>output_MAC_38_16, I17=>output_MAC_38_17, I18=>output_MAC_38_18, I19=>output_MAC_38_19, I20=>output_MAC_38_20, I21=>output_MAC_38_21, I22=>output_MAC_38_22, I23=>output_MAC_38_23, I24=>output_MAC_38_24, I25=>output_MAC_38_25, I26=>output_MAC_38_26, I27=>output_MAC_38_27, I28=>output_MAC_38_28, I29=>output_MAC_38_29, I30=>output_MAC_38_30, I31=>output_MAC_38_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_38);

	mux_row_39: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_39_0, I1=>output_MAC_39_1, I2=>output_MAC_39_2, I3=>output_MAC_39_3, I4=>output_MAC_39_4, I5=>output_MAC_39_5, I6=>output_MAC_39_6, I7=>output_MAC_39_7, I8=>output_MAC_39_8, I9=>output_MAC_39_9, I10=>output_MAC_39_10, I11=>output_MAC_39_11, I12=>output_MAC_39_12, I13=>output_MAC_39_13, I14=>output_MAC_39_14, I15=>output_MAC_39_15, I16=>output_MAC_39_16, I17=>output_MAC_39_17, I18=>output_MAC_39_18, I19=>output_MAC_39_19, I20=>output_MAC_39_20, I21=>output_MAC_39_21, I22=>output_MAC_39_22, I23=>output_MAC_39_23, I24=>output_MAC_39_24, I25=>output_MAC_39_25, I26=>output_MAC_39_26, I27=>output_MAC_39_27, I28=>output_MAC_39_28, I29=>output_MAC_39_29, I30=>output_MAC_39_30, I31=>output_MAC_39_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_39);

	mux_row_40: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_40_0, I1=>output_MAC_40_1, I2=>output_MAC_40_2, I3=>output_MAC_40_3, I4=>output_MAC_40_4, I5=>output_MAC_40_5, I6=>output_MAC_40_6, I7=>output_MAC_40_7, I8=>output_MAC_40_8, I9=>output_MAC_40_9, I10=>output_MAC_40_10, I11=>output_MAC_40_11, I12=>output_MAC_40_12, I13=>output_MAC_40_13, I14=>output_MAC_40_14, I15=>output_MAC_40_15, I16=>output_MAC_40_16, I17=>output_MAC_40_17, I18=>output_MAC_40_18, I19=>output_MAC_40_19, I20=>output_MAC_40_20, I21=>output_MAC_40_21, I22=>output_MAC_40_22, I23=>output_MAC_40_23, I24=>output_MAC_40_24, I25=>output_MAC_40_25, I26=>output_MAC_40_26, I27=>output_MAC_40_27, I28=>output_MAC_40_28, I29=>output_MAC_40_29, I30=>output_MAC_40_30, I31=>output_MAC_40_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_40);

	mux_row_41: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_41_0, I1=>output_MAC_41_1, I2=>output_MAC_41_2, I3=>output_MAC_41_3, I4=>output_MAC_41_4, I5=>output_MAC_41_5, I6=>output_MAC_41_6, I7=>output_MAC_41_7, I8=>output_MAC_41_8, I9=>output_MAC_41_9, I10=>output_MAC_41_10, I11=>output_MAC_41_11, I12=>output_MAC_41_12, I13=>output_MAC_41_13, I14=>output_MAC_41_14, I15=>output_MAC_41_15, I16=>output_MAC_41_16, I17=>output_MAC_41_17, I18=>output_MAC_41_18, I19=>output_MAC_41_19, I20=>output_MAC_41_20, I21=>output_MAC_41_21, I22=>output_MAC_41_22, I23=>output_MAC_41_23, I24=>output_MAC_41_24, I25=>output_MAC_41_25, I26=>output_MAC_41_26, I27=>output_MAC_41_27, I28=>output_MAC_41_28, I29=>output_MAC_41_29, I30=>output_MAC_41_30, I31=>output_MAC_41_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_41);

	mux_row_42: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_42_0, I1=>output_MAC_42_1, I2=>output_MAC_42_2, I3=>output_MAC_42_3, I4=>output_MAC_42_4, I5=>output_MAC_42_5, I6=>output_MAC_42_6, I7=>output_MAC_42_7, I8=>output_MAC_42_8, I9=>output_MAC_42_9, I10=>output_MAC_42_10, I11=>output_MAC_42_11, I12=>output_MAC_42_12, I13=>output_MAC_42_13, I14=>output_MAC_42_14, I15=>output_MAC_42_15, I16=>output_MAC_42_16, I17=>output_MAC_42_17, I18=>output_MAC_42_18, I19=>output_MAC_42_19, I20=>output_MAC_42_20, I21=>output_MAC_42_21, I22=>output_MAC_42_22, I23=>output_MAC_42_23, I24=>output_MAC_42_24, I25=>output_MAC_42_25, I26=>output_MAC_42_26, I27=>output_MAC_42_27, I28=>output_MAC_42_28, I29=>output_MAC_42_29, I30=>output_MAC_42_30, I31=>output_MAC_42_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_42);

	mux_row_43: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_43_0, I1=>output_MAC_43_1, I2=>output_MAC_43_2, I3=>output_MAC_43_3, I4=>output_MAC_43_4, I5=>output_MAC_43_5, I6=>output_MAC_43_6, I7=>output_MAC_43_7, I8=>output_MAC_43_8, I9=>output_MAC_43_9, I10=>output_MAC_43_10, I11=>output_MAC_43_11, I12=>output_MAC_43_12, I13=>output_MAC_43_13, I14=>output_MAC_43_14, I15=>output_MAC_43_15, I16=>output_MAC_43_16, I17=>output_MAC_43_17, I18=>output_MAC_43_18, I19=>output_MAC_43_19, I20=>output_MAC_43_20, I21=>output_MAC_43_21, I22=>output_MAC_43_22, I23=>output_MAC_43_23, I24=>output_MAC_43_24, I25=>output_MAC_43_25, I26=>output_MAC_43_26, I27=>output_MAC_43_27, I28=>output_MAC_43_28, I29=>output_MAC_43_29, I30=>output_MAC_43_30, I31=>output_MAC_43_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_43);

	mux_row_44: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_44_0, I1=>output_MAC_44_1, I2=>output_MAC_44_2, I3=>output_MAC_44_3, I4=>output_MAC_44_4, I5=>output_MAC_44_5, I6=>output_MAC_44_6, I7=>output_MAC_44_7, I8=>output_MAC_44_8, I9=>output_MAC_44_9, I10=>output_MAC_44_10, I11=>output_MAC_44_11, I12=>output_MAC_44_12, I13=>output_MAC_44_13, I14=>output_MAC_44_14, I15=>output_MAC_44_15, I16=>output_MAC_44_16, I17=>output_MAC_44_17, I18=>output_MAC_44_18, I19=>output_MAC_44_19, I20=>output_MAC_44_20, I21=>output_MAC_44_21, I22=>output_MAC_44_22, I23=>output_MAC_44_23, I24=>output_MAC_44_24, I25=>output_MAC_44_25, I26=>output_MAC_44_26, I27=>output_MAC_44_27, I28=>output_MAC_44_28, I29=>output_MAC_44_29, I30=>output_MAC_44_30, I31=>output_MAC_44_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_44);

	mux_row_45: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_45_0, I1=>output_MAC_45_1, I2=>output_MAC_45_2, I3=>output_MAC_45_3, I4=>output_MAC_45_4, I5=>output_MAC_45_5, I6=>output_MAC_45_6, I7=>output_MAC_45_7, I8=>output_MAC_45_8, I9=>output_MAC_45_9, I10=>output_MAC_45_10, I11=>output_MAC_45_11, I12=>output_MAC_45_12, I13=>output_MAC_45_13, I14=>output_MAC_45_14, I15=>output_MAC_45_15, I16=>output_MAC_45_16, I17=>output_MAC_45_17, I18=>output_MAC_45_18, I19=>output_MAC_45_19, I20=>output_MAC_45_20, I21=>output_MAC_45_21, I22=>output_MAC_45_22, I23=>output_MAC_45_23, I24=>output_MAC_45_24, I25=>output_MAC_45_25, I26=>output_MAC_45_26, I27=>output_MAC_45_27, I28=>output_MAC_45_28, I29=>output_MAC_45_29, I30=>output_MAC_45_30, I31=>output_MAC_45_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_45);

	mux_row_46: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_46_0, I1=>output_MAC_46_1, I2=>output_MAC_46_2, I3=>output_MAC_46_3, I4=>output_MAC_46_4, I5=>output_MAC_46_5, I6=>output_MAC_46_6, I7=>output_MAC_46_7, I8=>output_MAC_46_8, I9=>output_MAC_46_9, I10=>output_MAC_46_10, I11=>output_MAC_46_11, I12=>output_MAC_46_12, I13=>output_MAC_46_13, I14=>output_MAC_46_14, I15=>output_MAC_46_15, I16=>output_MAC_46_16, I17=>output_MAC_46_17, I18=>output_MAC_46_18, I19=>output_MAC_46_19, I20=>output_MAC_46_20, I21=>output_MAC_46_21, I22=>output_MAC_46_22, I23=>output_MAC_46_23, I24=>output_MAC_46_24, I25=>output_MAC_46_25, I26=>output_MAC_46_26, I27=>output_MAC_46_27, I28=>output_MAC_46_28, I29=>output_MAC_46_29, I30=>output_MAC_46_30, I31=>output_MAC_46_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_46);

	mux_row_47: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_47_0, I1=>output_MAC_47_1, I2=>output_MAC_47_2, I3=>output_MAC_47_3, I4=>output_MAC_47_4, I5=>output_MAC_47_5, I6=>output_MAC_47_6, I7=>output_MAC_47_7, I8=>output_MAC_47_8, I9=>output_MAC_47_9, I10=>output_MAC_47_10, I11=>output_MAC_47_11, I12=>output_MAC_47_12, I13=>output_MAC_47_13, I14=>output_MAC_47_14, I15=>output_MAC_47_15, I16=>output_MAC_47_16, I17=>output_MAC_47_17, I18=>output_MAC_47_18, I19=>output_MAC_47_19, I20=>output_MAC_47_20, I21=>output_MAC_47_21, I22=>output_MAC_47_22, I23=>output_MAC_47_23, I24=>output_MAC_47_24, I25=>output_MAC_47_25, I26=>output_MAC_47_26, I27=>output_MAC_47_27, I28=>output_MAC_47_28, I29=>output_MAC_47_29, I30=>output_MAC_47_30, I31=>output_MAC_47_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_47);

	mux_row_48: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_48_0, I1=>output_MAC_48_1, I2=>output_MAC_48_2, I3=>output_MAC_48_3, I4=>output_MAC_48_4, I5=>output_MAC_48_5, I6=>output_MAC_48_6, I7=>output_MAC_48_7, I8=>output_MAC_48_8, I9=>output_MAC_48_9, I10=>output_MAC_48_10, I11=>output_MAC_48_11, I12=>output_MAC_48_12, I13=>output_MAC_48_13, I14=>output_MAC_48_14, I15=>output_MAC_48_15, I16=>output_MAC_48_16, I17=>output_MAC_48_17, I18=>output_MAC_48_18, I19=>output_MAC_48_19, I20=>output_MAC_48_20, I21=>output_MAC_48_21, I22=>output_MAC_48_22, I23=>output_MAC_48_23, I24=>output_MAC_48_24, I25=>output_MAC_48_25, I26=>output_MAC_48_26, I27=>output_MAC_48_27, I28=>output_MAC_48_28, I29=>output_MAC_48_29, I30=>output_MAC_48_30, I31=>output_MAC_48_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_48);

	mux_row_49: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_49_0, I1=>output_MAC_49_1, I2=>output_MAC_49_2, I3=>output_MAC_49_3, I4=>output_MAC_49_4, I5=>output_MAC_49_5, I6=>output_MAC_49_6, I7=>output_MAC_49_7, I8=>output_MAC_49_8, I9=>output_MAC_49_9, I10=>output_MAC_49_10, I11=>output_MAC_49_11, I12=>output_MAC_49_12, I13=>output_MAC_49_13, I14=>output_MAC_49_14, I15=>output_MAC_49_15, I16=>output_MAC_49_16, I17=>output_MAC_49_17, I18=>output_MAC_49_18, I19=>output_MAC_49_19, I20=>output_MAC_49_20, I21=>output_MAC_49_21, I22=>output_MAC_49_22, I23=>output_MAC_49_23, I24=>output_MAC_49_24, I25=>output_MAC_49_25, I26=>output_MAC_49_26, I27=>output_MAC_49_27, I28=>output_MAC_49_28, I29=>output_MAC_49_29, I30=>output_MAC_49_30, I31=>output_MAC_49_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_49);

	mux_row_50: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_50_0, I1=>output_MAC_50_1, I2=>output_MAC_50_2, I3=>output_MAC_50_3, I4=>output_MAC_50_4, I5=>output_MAC_50_5, I6=>output_MAC_50_6, I7=>output_MAC_50_7, I8=>output_MAC_50_8, I9=>output_MAC_50_9, I10=>output_MAC_50_10, I11=>output_MAC_50_11, I12=>output_MAC_50_12, I13=>output_MAC_50_13, I14=>output_MAC_50_14, I15=>output_MAC_50_15, I16=>output_MAC_50_16, I17=>output_MAC_50_17, I18=>output_MAC_50_18, I19=>output_MAC_50_19, I20=>output_MAC_50_20, I21=>output_MAC_50_21, I22=>output_MAC_50_22, I23=>output_MAC_50_23, I24=>output_MAC_50_24, I25=>output_MAC_50_25, I26=>output_MAC_50_26, I27=>output_MAC_50_27, I28=>output_MAC_50_28, I29=>output_MAC_50_29, I30=>output_MAC_50_30, I31=>output_MAC_50_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_50);

	mux_row_51: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_51_0, I1=>output_MAC_51_1, I2=>output_MAC_51_2, I3=>output_MAC_51_3, I4=>output_MAC_51_4, I5=>output_MAC_51_5, I6=>output_MAC_51_6, I7=>output_MAC_51_7, I8=>output_MAC_51_8, I9=>output_MAC_51_9, I10=>output_MAC_51_10, I11=>output_MAC_51_11, I12=>output_MAC_51_12, I13=>output_MAC_51_13, I14=>output_MAC_51_14, I15=>output_MAC_51_15, I16=>output_MAC_51_16, I17=>output_MAC_51_17, I18=>output_MAC_51_18, I19=>output_MAC_51_19, I20=>output_MAC_51_20, I21=>output_MAC_51_21, I22=>output_MAC_51_22, I23=>output_MAC_51_23, I24=>output_MAC_51_24, I25=>output_MAC_51_25, I26=>output_MAC_51_26, I27=>output_MAC_51_27, I28=>output_MAC_51_28, I29=>output_MAC_51_29, I30=>output_MAC_51_30, I31=>output_MAC_51_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_51);

	mux_row_52: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_52_0, I1=>output_MAC_52_1, I2=>output_MAC_52_2, I3=>output_MAC_52_3, I4=>output_MAC_52_4, I5=>output_MAC_52_5, I6=>output_MAC_52_6, I7=>output_MAC_52_7, I8=>output_MAC_52_8, I9=>output_MAC_52_9, I10=>output_MAC_52_10, I11=>output_MAC_52_11, I12=>output_MAC_52_12, I13=>output_MAC_52_13, I14=>output_MAC_52_14, I15=>output_MAC_52_15, I16=>output_MAC_52_16, I17=>output_MAC_52_17, I18=>output_MAC_52_18, I19=>output_MAC_52_19, I20=>output_MAC_52_20, I21=>output_MAC_52_21, I22=>output_MAC_52_22, I23=>output_MAC_52_23, I24=>output_MAC_52_24, I25=>output_MAC_52_25, I26=>output_MAC_52_26, I27=>output_MAC_52_27, I28=>output_MAC_52_28, I29=>output_MAC_52_29, I30=>output_MAC_52_30, I31=>output_MAC_52_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_52);

	mux_row_53: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_53_0, I1=>output_MAC_53_1, I2=>output_MAC_53_2, I3=>output_MAC_53_3, I4=>output_MAC_53_4, I5=>output_MAC_53_5, I6=>output_MAC_53_6, I7=>output_MAC_53_7, I8=>output_MAC_53_8, I9=>output_MAC_53_9, I10=>output_MAC_53_10, I11=>output_MAC_53_11, I12=>output_MAC_53_12, I13=>output_MAC_53_13, I14=>output_MAC_53_14, I15=>output_MAC_53_15, I16=>output_MAC_53_16, I17=>output_MAC_53_17, I18=>output_MAC_53_18, I19=>output_MAC_53_19, I20=>output_MAC_53_20, I21=>output_MAC_53_21, I22=>output_MAC_53_22, I23=>output_MAC_53_23, I24=>output_MAC_53_24, I25=>output_MAC_53_25, I26=>output_MAC_53_26, I27=>output_MAC_53_27, I28=>output_MAC_53_28, I29=>output_MAC_53_29, I30=>output_MAC_53_30, I31=>output_MAC_53_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_53);

	mux_row_54: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_54_0, I1=>output_MAC_54_1, I2=>output_MAC_54_2, I3=>output_MAC_54_3, I4=>output_MAC_54_4, I5=>output_MAC_54_5, I6=>output_MAC_54_6, I7=>output_MAC_54_7, I8=>output_MAC_54_8, I9=>output_MAC_54_9, I10=>output_MAC_54_10, I11=>output_MAC_54_11, I12=>output_MAC_54_12, I13=>output_MAC_54_13, I14=>output_MAC_54_14, I15=>output_MAC_54_15, I16=>output_MAC_54_16, I17=>output_MAC_54_17, I18=>output_MAC_54_18, I19=>output_MAC_54_19, I20=>output_MAC_54_20, I21=>output_MAC_54_21, I22=>output_MAC_54_22, I23=>output_MAC_54_23, I24=>output_MAC_54_24, I25=>output_MAC_54_25, I26=>output_MAC_54_26, I27=>output_MAC_54_27, I28=>output_MAC_54_28, I29=>output_MAC_54_29, I30=>output_MAC_54_30, I31=>output_MAC_54_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_54);

	mux_row_55: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_55_0, I1=>output_MAC_55_1, I2=>output_MAC_55_2, I3=>output_MAC_55_3, I4=>output_MAC_55_4, I5=>output_MAC_55_5, I6=>output_MAC_55_6, I7=>output_MAC_55_7, I8=>output_MAC_55_8, I9=>output_MAC_55_9, I10=>output_MAC_55_10, I11=>output_MAC_55_11, I12=>output_MAC_55_12, I13=>output_MAC_55_13, I14=>output_MAC_55_14, I15=>output_MAC_55_15, I16=>output_MAC_55_16, I17=>output_MAC_55_17, I18=>output_MAC_55_18, I19=>output_MAC_55_19, I20=>output_MAC_55_20, I21=>output_MAC_55_21, I22=>output_MAC_55_22, I23=>output_MAC_55_23, I24=>output_MAC_55_24, I25=>output_MAC_55_25, I26=>output_MAC_55_26, I27=>output_MAC_55_27, I28=>output_MAC_55_28, I29=>output_MAC_55_29, I30=>output_MAC_55_30, I31=>output_MAC_55_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_55);

	mux_row_56: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_56_0, I1=>output_MAC_56_1, I2=>output_MAC_56_2, I3=>output_MAC_56_3, I4=>output_MAC_56_4, I5=>output_MAC_56_5, I6=>output_MAC_56_6, I7=>output_MAC_56_7, I8=>output_MAC_56_8, I9=>output_MAC_56_9, I10=>output_MAC_56_10, I11=>output_MAC_56_11, I12=>output_MAC_56_12, I13=>output_MAC_56_13, I14=>output_MAC_56_14, I15=>output_MAC_56_15, I16=>output_MAC_56_16, I17=>output_MAC_56_17, I18=>output_MAC_56_18, I19=>output_MAC_56_19, I20=>output_MAC_56_20, I21=>output_MAC_56_21, I22=>output_MAC_56_22, I23=>output_MAC_56_23, I24=>output_MAC_56_24, I25=>output_MAC_56_25, I26=>output_MAC_56_26, I27=>output_MAC_56_27, I28=>output_MAC_56_28, I29=>output_MAC_56_29, I30=>output_MAC_56_30, I31=>output_MAC_56_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_56);

	mux_row_57: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_57_0, I1=>output_MAC_57_1, I2=>output_MAC_57_2, I3=>output_MAC_57_3, I4=>output_MAC_57_4, I5=>output_MAC_57_5, I6=>output_MAC_57_6, I7=>output_MAC_57_7, I8=>output_MAC_57_8, I9=>output_MAC_57_9, I10=>output_MAC_57_10, I11=>output_MAC_57_11, I12=>output_MAC_57_12, I13=>output_MAC_57_13, I14=>output_MAC_57_14, I15=>output_MAC_57_15, I16=>output_MAC_57_16, I17=>output_MAC_57_17, I18=>output_MAC_57_18, I19=>output_MAC_57_19, I20=>output_MAC_57_20, I21=>output_MAC_57_21, I22=>output_MAC_57_22, I23=>output_MAC_57_23, I24=>output_MAC_57_24, I25=>output_MAC_57_25, I26=>output_MAC_57_26, I27=>output_MAC_57_27, I28=>output_MAC_57_28, I29=>output_MAC_57_29, I30=>output_MAC_57_30, I31=>output_MAC_57_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_57);

	mux_row_58: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_58_0, I1=>output_MAC_58_1, I2=>output_MAC_58_2, I3=>output_MAC_58_3, I4=>output_MAC_58_4, I5=>output_MAC_58_5, I6=>output_MAC_58_6, I7=>output_MAC_58_7, I8=>output_MAC_58_8, I9=>output_MAC_58_9, I10=>output_MAC_58_10, I11=>output_MAC_58_11, I12=>output_MAC_58_12, I13=>output_MAC_58_13, I14=>output_MAC_58_14, I15=>output_MAC_58_15, I16=>output_MAC_58_16, I17=>output_MAC_58_17, I18=>output_MAC_58_18, I19=>output_MAC_58_19, I20=>output_MAC_58_20, I21=>output_MAC_58_21, I22=>output_MAC_58_22, I23=>output_MAC_58_23, I24=>output_MAC_58_24, I25=>output_MAC_58_25, I26=>output_MAC_58_26, I27=>output_MAC_58_27, I28=>output_MAC_58_28, I29=>output_MAC_58_29, I30=>output_MAC_58_30, I31=>output_MAC_58_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_58);

	mux_row_59: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_59_0, I1=>output_MAC_59_1, I2=>output_MAC_59_2, I3=>output_MAC_59_3, I4=>output_MAC_59_4, I5=>output_MAC_59_5, I6=>output_MAC_59_6, I7=>output_MAC_59_7, I8=>output_MAC_59_8, I9=>output_MAC_59_9, I10=>output_MAC_59_10, I11=>output_MAC_59_11, I12=>output_MAC_59_12, I13=>output_MAC_59_13, I14=>output_MAC_59_14, I15=>output_MAC_59_15, I16=>output_MAC_59_16, I17=>output_MAC_59_17, I18=>output_MAC_59_18, I19=>output_MAC_59_19, I20=>output_MAC_59_20, I21=>output_MAC_59_21, I22=>output_MAC_59_22, I23=>output_MAC_59_23, I24=>output_MAC_59_24, I25=>output_MAC_59_25, I26=>output_MAC_59_26, I27=>output_MAC_59_27, I28=>output_MAC_59_28, I29=>output_MAC_59_29, I30=>output_MAC_59_30, I31=>output_MAC_59_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_59);

	mux_row_60: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_60_0, I1=>output_MAC_60_1, I2=>output_MAC_60_2, I3=>output_MAC_60_3, I4=>output_MAC_60_4, I5=>output_MAC_60_5, I6=>output_MAC_60_6, I7=>output_MAC_60_7, I8=>output_MAC_60_8, I9=>output_MAC_60_9, I10=>output_MAC_60_10, I11=>output_MAC_60_11, I12=>output_MAC_60_12, I13=>output_MAC_60_13, I14=>output_MAC_60_14, I15=>output_MAC_60_15, I16=>output_MAC_60_16, I17=>output_MAC_60_17, I18=>output_MAC_60_18, I19=>output_MAC_60_19, I20=>output_MAC_60_20, I21=>output_MAC_60_21, I22=>output_MAC_60_22, I23=>output_MAC_60_23, I24=>output_MAC_60_24, I25=>output_MAC_60_25, I26=>output_MAC_60_26, I27=>output_MAC_60_27, I28=>output_MAC_60_28, I29=>output_MAC_60_29, I30=>output_MAC_60_30, I31=>output_MAC_60_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_60);

	mux_row_61: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_61_0, I1=>output_MAC_61_1, I2=>output_MAC_61_2, I3=>output_MAC_61_3, I4=>output_MAC_61_4, I5=>output_MAC_61_5, I6=>output_MAC_61_6, I7=>output_MAC_61_7, I8=>output_MAC_61_8, I9=>output_MAC_61_9, I10=>output_MAC_61_10, I11=>output_MAC_61_11, I12=>output_MAC_61_12, I13=>output_MAC_61_13, I14=>output_MAC_61_14, I15=>output_MAC_61_15, I16=>output_MAC_61_16, I17=>output_MAC_61_17, I18=>output_MAC_61_18, I19=>output_MAC_61_19, I20=>output_MAC_61_20, I21=>output_MAC_61_21, I22=>output_MAC_61_22, I23=>output_MAC_61_23, I24=>output_MAC_61_24, I25=>output_MAC_61_25, I26=>output_MAC_61_26, I27=>output_MAC_61_27, I28=>output_MAC_61_28, I29=>output_MAC_61_29, I30=>output_MAC_61_30, I31=>output_MAC_61_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_61);

	mux_row_62: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_62_0, I1=>output_MAC_62_1, I2=>output_MAC_62_2, I3=>output_MAC_62_3, I4=>output_MAC_62_4, I5=>output_MAC_62_5, I6=>output_MAC_62_6, I7=>output_MAC_62_7, I8=>output_MAC_62_8, I9=>output_MAC_62_9, I10=>output_MAC_62_10, I11=>output_MAC_62_11, I12=>output_MAC_62_12, I13=>output_MAC_62_13, I14=>output_MAC_62_14, I15=>output_MAC_62_15, I16=>output_MAC_62_16, I17=>output_MAC_62_17, I18=>output_MAC_62_18, I19=>output_MAC_62_19, I20=>output_MAC_62_20, I21=>output_MAC_62_21, I22=>output_MAC_62_22, I23=>output_MAC_62_23, I24=>output_MAC_62_24, I25=>output_MAC_62_25, I26=>output_MAC_62_26, I27=>output_MAC_62_27, I28=>output_MAC_62_28, I29=>output_MAC_62_29, I30=>output_MAC_62_30, I31=>output_MAC_62_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_62);

	mux_row_63: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_63_0, I1=>output_MAC_63_1, I2=>output_MAC_63_2, I3=>output_MAC_63_3, I4=>output_MAC_63_4, I5=>output_MAC_63_5, I6=>output_MAC_63_6, I7=>output_MAC_63_7, I8=>output_MAC_63_8, I9=>output_MAC_63_9, I10=>output_MAC_63_10, I11=>output_MAC_63_11, I12=>output_MAC_63_12, I13=>output_MAC_63_13, I14=>output_MAC_63_14, I15=>output_MAC_63_15, I16=>output_MAC_63_16, I17=>output_MAC_63_17, I18=>output_MAC_63_18, I19=>output_MAC_63_19, I20=>output_MAC_63_20, I21=>output_MAC_63_21, I22=>output_MAC_63_22, I23=>output_MAC_63_23, I24=>output_MAC_63_24, I25=>output_MAC_63_25, I26=>output_MAC_63_26, I27=>output_MAC_63_27, I28=>output_MAC_63_28, I29=>output_MAC_63_29, I30=>output_MAC_63_30, I31=>output_MAC_63_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_63);

	mux_row_64: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_64_0, I1=>output_MAC_64_1, I2=>output_MAC_64_2, I3=>output_MAC_64_3, I4=>output_MAC_64_4, I5=>output_MAC_64_5, I6=>output_MAC_64_6, I7=>output_MAC_64_7, I8=>output_MAC_64_8, I9=>output_MAC_64_9, I10=>output_MAC_64_10, I11=>output_MAC_64_11, I12=>output_MAC_64_12, I13=>output_MAC_64_13, I14=>output_MAC_64_14, I15=>output_MAC_64_15, I16=>output_MAC_64_16, I17=>output_MAC_64_17, I18=>output_MAC_64_18, I19=>output_MAC_64_19, I20=>output_MAC_64_20, I21=>output_MAC_64_21, I22=>output_MAC_64_22, I23=>output_MAC_64_23, I24=>output_MAC_64_24, I25=>output_MAC_64_25, I26=>output_MAC_64_26, I27=>output_MAC_64_27, I28=>output_MAC_64_28, I29=>output_MAC_64_29, I30=>output_MAC_64_30, I31=>output_MAC_64_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_64);

	mux_row_65: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_65_0, I1=>output_MAC_65_1, I2=>output_MAC_65_2, I3=>output_MAC_65_3, I4=>output_MAC_65_4, I5=>output_MAC_65_5, I6=>output_MAC_65_6, I7=>output_MAC_65_7, I8=>output_MAC_65_8, I9=>output_MAC_65_9, I10=>output_MAC_65_10, I11=>output_MAC_65_11, I12=>output_MAC_65_12, I13=>output_MAC_65_13, I14=>output_MAC_65_14, I15=>output_MAC_65_15, I16=>output_MAC_65_16, I17=>output_MAC_65_17, I18=>output_MAC_65_18, I19=>output_MAC_65_19, I20=>output_MAC_65_20, I21=>output_MAC_65_21, I22=>output_MAC_65_22, I23=>output_MAC_65_23, I24=>output_MAC_65_24, I25=>output_MAC_65_25, I26=>output_MAC_65_26, I27=>output_MAC_65_27, I28=>output_MAC_65_28, I29=>output_MAC_65_29, I30=>output_MAC_65_30, I31=>output_MAC_65_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_65);

	mux_row_66: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_66_0, I1=>output_MAC_66_1, I2=>output_MAC_66_2, I3=>output_MAC_66_3, I4=>output_MAC_66_4, I5=>output_MAC_66_5, I6=>output_MAC_66_6, I7=>output_MAC_66_7, I8=>output_MAC_66_8, I9=>output_MAC_66_9, I10=>output_MAC_66_10, I11=>output_MAC_66_11, I12=>output_MAC_66_12, I13=>output_MAC_66_13, I14=>output_MAC_66_14, I15=>output_MAC_66_15, I16=>output_MAC_66_16, I17=>output_MAC_66_17, I18=>output_MAC_66_18, I19=>output_MAC_66_19, I20=>output_MAC_66_20, I21=>output_MAC_66_21, I22=>output_MAC_66_22, I23=>output_MAC_66_23, I24=>output_MAC_66_24, I25=>output_MAC_66_25, I26=>output_MAC_66_26, I27=>output_MAC_66_27, I28=>output_MAC_66_28, I29=>output_MAC_66_29, I30=>output_MAC_66_30, I31=>output_MAC_66_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_66);

	mux_row_67: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_67_0, I1=>output_MAC_67_1, I2=>output_MAC_67_2, I3=>output_MAC_67_3, I4=>output_MAC_67_4, I5=>output_MAC_67_5, I6=>output_MAC_67_6, I7=>output_MAC_67_7, I8=>output_MAC_67_8, I9=>output_MAC_67_9, I10=>output_MAC_67_10, I11=>output_MAC_67_11, I12=>output_MAC_67_12, I13=>output_MAC_67_13, I14=>output_MAC_67_14, I15=>output_MAC_67_15, I16=>output_MAC_67_16, I17=>output_MAC_67_17, I18=>output_MAC_67_18, I19=>output_MAC_67_19, I20=>output_MAC_67_20, I21=>output_MAC_67_21, I22=>output_MAC_67_22, I23=>output_MAC_67_23, I24=>output_MAC_67_24, I25=>output_MAC_67_25, I26=>output_MAC_67_26, I27=>output_MAC_67_27, I28=>output_MAC_67_28, I29=>output_MAC_67_29, I30=>output_MAC_67_30, I31=>output_MAC_67_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_67);

	mux_row_68: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_68_0, I1=>output_MAC_68_1, I2=>output_MAC_68_2, I3=>output_MAC_68_3, I4=>output_MAC_68_4, I5=>output_MAC_68_5, I6=>output_MAC_68_6, I7=>output_MAC_68_7, I8=>output_MAC_68_8, I9=>output_MAC_68_9, I10=>output_MAC_68_10, I11=>output_MAC_68_11, I12=>output_MAC_68_12, I13=>output_MAC_68_13, I14=>output_MAC_68_14, I15=>output_MAC_68_15, I16=>output_MAC_68_16, I17=>output_MAC_68_17, I18=>output_MAC_68_18, I19=>output_MAC_68_19, I20=>output_MAC_68_20, I21=>output_MAC_68_21, I22=>output_MAC_68_22, I23=>output_MAC_68_23, I24=>output_MAC_68_24, I25=>output_MAC_68_25, I26=>output_MAC_68_26, I27=>output_MAC_68_27, I28=>output_MAC_68_28, I29=>output_MAC_68_29, I30=>output_MAC_68_30, I31=>output_MAC_68_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_68);

	mux_row_69: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_69_0, I1=>output_MAC_69_1, I2=>output_MAC_69_2, I3=>output_MAC_69_3, I4=>output_MAC_69_4, I5=>output_MAC_69_5, I6=>output_MAC_69_6, I7=>output_MAC_69_7, I8=>output_MAC_69_8, I9=>output_MAC_69_9, I10=>output_MAC_69_10, I11=>output_MAC_69_11, I12=>output_MAC_69_12, I13=>output_MAC_69_13, I14=>output_MAC_69_14, I15=>output_MAC_69_15, I16=>output_MAC_69_16, I17=>output_MAC_69_17, I18=>output_MAC_69_18, I19=>output_MAC_69_19, I20=>output_MAC_69_20, I21=>output_MAC_69_21, I22=>output_MAC_69_22, I23=>output_MAC_69_23, I24=>output_MAC_69_24, I25=>output_MAC_69_25, I26=>output_MAC_69_26, I27=>output_MAC_69_27, I28=>output_MAC_69_28, I29=>output_MAC_69_29, I30=>output_MAC_69_30, I31=>output_MAC_69_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_69);

	mux_row_70: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_70_0, I1=>output_MAC_70_1, I2=>output_MAC_70_2, I3=>output_MAC_70_3, I4=>output_MAC_70_4, I5=>output_MAC_70_5, I6=>output_MAC_70_6, I7=>output_MAC_70_7, I8=>output_MAC_70_8, I9=>output_MAC_70_9, I10=>output_MAC_70_10, I11=>output_MAC_70_11, I12=>output_MAC_70_12, I13=>output_MAC_70_13, I14=>output_MAC_70_14, I15=>output_MAC_70_15, I16=>output_MAC_70_16, I17=>output_MAC_70_17, I18=>output_MAC_70_18, I19=>output_MAC_70_19, I20=>output_MAC_70_20, I21=>output_MAC_70_21, I22=>output_MAC_70_22, I23=>output_MAC_70_23, I24=>output_MAC_70_24, I25=>output_MAC_70_25, I26=>output_MAC_70_26, I27=>output_MAC_70_27, I28=>output_MAC_70_28, I29=>output_MAC_70_29, I30=>output_MAC_70_30, I31=>output_MAC_70_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_70);

	mux_row_71: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_71_0, I1=>output_MAC_71_1, I2=>output_MAC_71_2, I3=>output_MAC_71_3, I4=>output_MAC_71_4, I5=>output_MAC_71_5, I6=>output_MAC_71_6, I7=>output_MAC_71_7, I8=>output_MAC_71_8, I9=>output_MAC_71_9, I10=>output_MAC_71_10, I11=>output_MAC_71_11, I12=>output_MAC_71_12, I13=>output_MAC_71_13, I14=>output_MAC_71_14, I15=>output_MAC_71_15, I16=>output_MAC_71_16, I17=>output_MAC_71_17, I18=>output_MAC_71_18, I19=>output_MAC_71_19, I20=>output_MAC_71_20, I21=>output_MAC_71_21, I22=>output_MAC_71_22, I23=>output_MAC_71_23, I24=>output_MAC_71_24, I25=>output_MAC_71_25, I26=>output_MAC_71_26, I27=>output_MAC_71_27, I28=>output_MAC_71_28, I29=>output_MAC_71_29, I30=>output_MAC_71_30, I31=>output_MAC_71_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_71);

	mux_row_72: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_72_0, I1=>output_MAC_72_1, I2=>output_MAC_72_2, I3=>output_MAC_72_3, I4=>output_MAC_72_4, I5=>output_MAC_72_5, I6=>output_MAC_72_6, I7=>output_MAC_72_7, I8=>output_MAC_72_8, I9=>output_MAC_72_9, I10=>output_MAC_72_10, I11=>output_MAC_72_11, I12=>output_MAC_72_12, I13=>output_MAC_72_13, I14=>output_MAC_72_14, I15=>output_MAC_72_15, I16=>output_MAC_72_16, I17=>output_MAC_72_17, I18=>output_MAC_72_18, I19=>output_MAC_72_19, I20=>output_MAC_72_20, I21=>output_MAC_72_21, I22=>output_MAC_72_22, I23=>output_MAC_72_23, I24=>output_MAC_72_24, I25=>output_MAC_72_25, I26=>output_MAC_72_26, I27=>output_MAC_72_27, I28=>output_MAC_72_28, I29=>output_MAC_72_29, I30=>output_MAC_72_30, I31=>output_MAC_72_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_72);

	mux_row_73: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_73_0, I1=>output_MAC_73_1, I2=>output_MAC_73_2, I3=>output_MAC_73_3, I4=>output_MAC_73_4, I5=>output_MAC_73_5, I6=>output_MAC_73_6, I7=>output_MAC_73_7, I8=>output_MAC_73_8, I9=>output_MAC_73_9, I10=>output_MAC_73_10, I11=>output_MAC_73_11, I12=>output_MAC_73_12, I13=>output_MAC_73_13, I14=>output_MAC_73_14, I15=>output_MAC_73_15, I16=>output_MAC_73_16, I17=>output_MAC_73_17, I18=>output_MAC_73_18, I19=>output_MAC_73_19, I20=>output_MAC_73_20, I21=>output_MAC_73_21, I22=>output_MAC_73_22, I23=>output_MAC_73_23, I24=>output_MAC_73_24, I25=>output_MAC_73_25, I26=>output_MAC_73_26, I27=>output_MAC_73_27, I28=>output_MAC_73_28, I29=>output_MAC_73_29, I30=>output_MAC_73_30, I31=>output_MAC_73_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_73);

	mux_row_74: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_74_0, I1=>output_MAC_74_1, I2=>output_MAC_74_2, I3=>output_MAC_74_3, I4=>output_MAC_74_4, I5=>output_MAC_74_5, I6=>output_MAC_74_6, I7=>output_MAC_74_7, I8=>output_MAC_74_8, I9=>output_MAC_74_9, I10=>output_MAC_74_10, I11=>output_MAC_74_11, I12=>output_MAC_74_12, I13=>output_MAC_74_13, I14=>output_MAC_74_14, I15=>output_MAC_74_15, I16=>output_MAC_74_16, I17=>output_MAC_74_17, I18=>output_MAC_74_18, I19=>output_MAC_74_19, I20=>output_MAC_74_20, I21=>output_MAC_74_21, I22=>output_MAC_74_22, I23=>output_MAC_74_23, I24=>output_MAC_74_24, I25=>output_MAC_74_25, I26=>output_MAC_74_26, I27=>output_MAC_74_27, I28=>output_MAC_74_28, I29=>output_MAC_74_29, I30=>output_MAC_74_30, I31=>output_MAC_74_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_74);

	mux_row_75: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_75_0, I1=>output_MAC_75_1, I2=>output_MAC_75_2, I3=>output_MAC_75_3, I4=>output_MAC_75_4, I5=>output_MAC_75_5, I6=>output_MAC_75_6, I7=>output_MAC_75_7, I8=>output_MAC_75_8, I9=>output_MAC_75_9, I10=>output_MAC_75_10, I11=>output_MAC_75_11, I12=>output_MAC_75_12, I13=>output_MAC_75_13, I14=>output_MAC_75_14, I15=>output_MAC_75_15, I16=>output_MAC_75_16, I17=>output_MAC_75_17, I18=>output_MAC_75_18, I19=>output_MAC_75_19, I20=>output_MAC_75_20, I21=>output_MAC_75_21, I22=>output_MAC_75_22, I23=>output_MAC_75_23, I24=>output_MAC_75_24, I25=>output_MAC_75_25, I26=>output_MAC_75_26, I27=>output_MAC_75_27, I28=>output_MAC_75_28, I29=>output_MAC_75_29, I30=>output_MAC_75_30, I31=>output_MAC_75_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_75);

	mux_row_76: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_76_0, I1=>output_MAC_76_1, I2=>output_MAC_76_2, I3=>output_MAC_76_3, I4=>output_MAC_76_4, I5=>output_MAC_76_5, I6=>output_MAC_76_6, I7=>output_MAC_76_7, I8=>output_MAC_76_8, I9=>output_MAC_76_9, I10=>output_MAC_76_10, I11=>output_MAC_76_11, I12=>output_MAC_76_12, I13=>output_MAC_76_13, I14=>output_MAC_76_14, I15=>output_MAC_76_15, I16=>output_MAC_76_16, I17=>output_MAC_76_17, I18=>output_MAC_76_18, I19=>output_MAC_76_19, I20=>output_MAC_76_20, I21=>output_MAC_76_21, I22=>output_MAC_76_22, I23=>output_MAC_76_23, I24=>output_MAC_76_24, I25=>output_MAC_76_25, I26=>output_MAC_76_26, I27=>output_MAC_76_27, I28=>output_MAC_76_28, I29=>output_MAC_76_29, I30=>output_MAC_76_30, I31=>output_MAC_76_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_76);

	mux_row_77: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_77_0, I1=>output_MAC_77_1, I2=>output_MAC_77_2, I3=>output_MAC_77_3, I4=>output_MAC_77_4, I5=>output_MAC_77_5, I6=>output_MAC_77_6, I7=>output_MAC_77_7, I8=>output_MAC_77_8, I9=>output_MAC_77_9, I10=>output_MAC_77_10, I11=>output_MAC_77_11, I12=>output_MAC_77_12, I13=>output_MAC_77_13, I14=>output_MAC_77_14, I15=>output_MAC_77_15, I16=>output_MAC_77_16, I17=>output_MAC_77_17, I18=>output_MAC_77_18, I19=>output_MAC_77_19, I20=>output_MAC_77_20, I21=>output_MAC_77_21, I22=>output_MAC_77_22, I23=>output_MAC_77_23, I24=>output_MAC_77_24, I25=>output_MAC_77_25, I26=>output_MAC_77_26, I27=>output_MAC_77_27, I28=>output_MAC_77_28, I29=>output_MAC_77_29, I30=>output_MAC_77_30, I31=>output_MAC_77_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_77);

	mux_row_78: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_78_0, I1=>output_MAC_78_1, I2=>output_MAC_78_2, I3=>output_MAC_78_3, I4=>output_MAC_78_4, I5=>output_MAC_78_5, I6=>output_MAC_78_6, I7=>output_MAC_78_7, I8=>output_MAC_78_8, I9=>output_MAC_78_9, I10=>output_MAC_78_10, I11=>output_MAC_78_11, I12=>output_MAC_78_12, I13=>output_MAC_78_13, I14=>output_MAC_78_14, I15=>output_MAC_78_15, I16=>output_MAC_78_16, I17=>output_MAC_78_17, I18=>output_MAC_78_18, I19=>output_MAC_78_19, I20=>output_MAC_78_20, I21=>output_MAC_78_21, I22=>output_MAC_78_22, I23=>output_MAC_78_23, I24=>output_MAC_78_24, I25=>output_MAC_78_25, I26=>output_MAC_78_26, I27=>output_MAC_78_27, I28=>output_MAC_78_28, I29=>output_MAC_78_29, I30=>output_MAC_78_30, I31=>output_MAC_78_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_78);

	mux_row_79: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_79_0, I1=>output_MAC_79_1, I2=>output_MAC_79_2, I3=>output_MAC_79_3, I4=>output_MAC_79_4, I5=>output_MAC_79_5, I6=>output_MAC_79_6, I7=>output_MAC_79_7, I8=>output_MAC_79_8, I9=>output_MAC_79_9, I10=>output_MAC_79_10, I11=>output_MAC_79_11, I12=>output_MAC_79_12, I13=>output_MAC_79_13, I14=>output_MAC_79_14, I15=>output_MAC_79_15, I16=>output_MAC_79_16, I17=>output_MAC_79_17, I18=>output_MAC_79_18, I19=>output_MAC_79_19, I20=>output_MAC_79_20, I21=>output_MAC_79_21, I22=>output_MAC_79_22, I23=>output_MAC_79_23, I24=>output_MAC_79_24, I25=>output_MAC_79_25, I26=>output_MAC_79_26, I27=>output_MAC_79_27, I28=>output_MAC_79_28, I29=>output_MAC_79_29, I30=>output_MAC_79_30, I31=>output_MAC_79_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_79);

	mux_row_80: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_80_0, I1=>output_MAC_80_1, I2=>output_MAC_80_2, I3=>output_MAC_80_3, I4=>output_MAC_80_4, I5=>output_MAC_80_5, I6=>output_MAC_80_6, I7=>output_MAC_80_7, I8=>output_MAC_80_8, I9=>output_MAC_80_9, I10=>output_MAC_80_10, I11=>output_MAC_80_11, I12=>output_MAC_80_12, I13=>output_MAC_80_13, I14=>output_MAC_80_14, I15=>output_MAC_80_15, I16=>output_MAC_80_16, I17=>output_MAC_80_17, I18=>output_MAC_80_18, I19=>output_MAC_80_19, I20=>output_MAC_80_20, I21=>output_MAC_80_21, I22=>output_MAC_80_22, I23=>output_MAC_80_23, I24=>output_MAC_80_24, I25=>output_MAC_80_25, I26=>output_MAC_80_26, I27=>output_MAC_80_27, I28=>output_MAC_80_28, I29=>output_MAC_80_29, I30=>output_MAC_80_30, I31=>output_MAC_80_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_80);

	mux_row_81: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_81_0, I1=>output_MAC_81_1, I2=>output_MAC_81_2, I3=>output_MAC_81_3, I4=>output_MAC_81_4, I5=>output_MAC_81_5, I6=>output_MAC_81_6, I7=>output_MAC_81_7, I8=>output_MAC_81_8, I9=>output_MAC_81_9, I10=>output_MAC_81_10, I11=>output_MAC_81_11, I12=>output_MAC_81_12, I13=>output_MAC_81_13, I14=>output_MAC_81_14, I15=>output_MAC_81_15, I16=>output_MAC_81_16, I17=>output_MAC_81_17, I18=>output_MAC_81_18, I19=>output_MAC_81_19, I20=>output_MAC_81_20, I21=>output_MAC_81_21, I22=>output_MAC_81_22, I23=>output_MAC_81_23, I24=>output_MAC_81_24, I25=>output_MAC_81_25, I26=>output_MAC_81_26, I27=>output_MAC_81_27, I28=>output_MAC_81_28, I29=>output_MAC_81_29, I30=>output_MAC_81_30, I31=>output_MAC_81_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_81);

	mux_row_82: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_82_0, I1=>output_MAC_82_1, I2=>output_MAC_82_2, I3=>output_MAC_82_3, I4=>output_MAC_82_4, I5=>output_MAC_82_5, I6=>output_MAC_82_6, I7=>output_MAC_82_7, I8=>output_MAC_82_8, I9=>output_MAC_82_9, I10=>output_MAC_82_10, I11=>output_MAC_82_11, I12=>output_MAC_82_12, I13=>output_MAC_82_13, I14=>output_MAC_82_14, I15=>output_MAC_82_15, I16=>output_MAC_82_16, I17=>output_MAC_82_17, I18=>output_MAC_82_18, I19=>output_MAC_82_19, I20=>output_MAC_82_20, I21=>output_MAC_82_21, I22=>output_MAC_82_22, I23=>output_MAC_82_23, I24=>output_MAC_82_24, I25=>output_MAC_82_25, I26=>output_MAC_82_26, I27=>output_MAC_82_27, I28=>output_MAC_82_28, I29=>output_MAC_82_29, I30=>output_MAC_82_30, I31=>output_MAC_82_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_82);

	mux_row_83: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_83_0, I1=>output_MAC_83_1, I2=>output_MAC_83_2, I3=>output_MAC_83_3, I4=>output_MAC_83_4, I5=>output_MAC_83_5, I6=>output_MAC_83_6, I7=>output_MAC_83_7, I8=>output_MAC_83_8, I9=>output_MAC_83_9, I10=>output_MAC_83_10, I11=>output_MAC_83_11, I12=>output_MAC_83_12, I13=>output_MAC_83_13, I14=>output_MAC_83_14, I15=>output_MAC_83_15, I16=>output_MAC_83_16, I17=>output_MAC_83_17, I18=>output_MAC_83_18, I19=>output_MAC_83_19, I20=>output_MAC_83_20, I21=>output_MAC_83_21, I22=>output_MAC_83_22, I23=>output_MAC_83_23, I24=>output_MAC_83_24, I25=>output_MAC_83_25, I26=>output_MAC_83_26, I27=>output_MAC_83_27, I28=>output_MAC_83_28, I29=>output_MAC_83_29, I30=>output_MAC_83_30, I31=>output_MAC_83_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_83);

	mux_row_84: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_84_0, I1=>output_MAC_84_1, I2=>output_MAC_84_2, I3=>output_MAC_84_3, I4=>output_MAC_84_4, I5=>output_MAC_84_5, I6=>output_MAC_84_6, I7=>output_MAC_84_7, I8=>output_MAC_84_8, I9=>output_MAC_84_9, I10=>output_MAC_84_10, I11=>output_MAC_84_11, I12=>output_MAC_84_12, I13=>output_MAC_84_13, I14=>output_MAC_84_14, I15=>output_MAC_84_15, I16=>output_MAC_84_16, I17=>output_MAC_84_17, I18=>output_MAC_84_18, I19=>output_MAC_84_19, I20=>output_MAC_84_20, I21=>output_MAC_84_21, I22=>output_MAC_84_22, I23=>output_MAC_84_23, I24=>output_MAC_84_24, I25=>output_MAC_84_25, I26=>output_MAC_84_26, I27=>output_MAC_84_27, I28=>output_MAC_84_28, I29=>output_MAC_84_29, I30=>output_MAC_84_30, I31=>output_MAC_84_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_84);

	mux_row_85: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_85_0, I1=>output_MAC_85_1, I2=>output_MAC_85_2, I3=>output_MAC_85_3, I4=>output_MAC_85_4, I5=>output_MAC_85_5, I6=>output_MAC_85_6, I7=>output_MAC_85_7, I8=>output_MAC_85_8, I9=>output_MAC_85_9, I10=>output_MAC_85_10, I11=>output_MAC_85_11, I12=>output_MAC_85_12, I13=>output_MAC_85_13, I14=>output_MAC_85_14, I15=>output_MAC_85_15, I16=>output_MAC_85_16, I17=>output_MAC_85_17, I18=>output_MAC_85_18, I19=>output_MAC_85_19, I20=>output_MAC_85_20, I21=>output_MAC_85_21, I22=>output_MAC_85_22, I23=>output_MAC_85_23, I24=>output_MAC_85_24, I25=>output_MAC_85_25, I26=>output_MAC_85_26, I27=>output_MAC_85_27, I28=>output_MAC_85_28, I29=>output_MAC_85_29, I30=>output_MAC_85_30, I31=>output_MAC_85_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_85);

	mux_row_86: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_86_0, I1=>output_MAC_86_1, I2=>output_MAC_86_2, I3=>output_MAC_86_3, I4=>output_MAC_86_4, I5=>output_MAC_86_5, I6=>output_MAC_86_6, I7=>output_MAC_86_7, I8=>output_MAC_86_8, I9=>output_MAC_86_9, I10=>output_MAC_86_10, I11=>output_MAC_86_11, I12=>output_MAC_86_12, I13=>output_MAC_86_13, I14=>output_MAC_86_14, I15=>output_MAC_86_15, I16=>output_MAC_86_16, I17=>output_MAC_86_17, I18=>output_MAC_86_18, I19=>output_MAC_86_19, I20=>output_MAC_86_20, I21=>output_MAC_86_21, I22=>output_MAC_86_22, I23=>output_MAC_86_23, I24=>output_MAC_86_24, I25=>output_MAC_86_25, I26=>output_MAC_86_26, I27=>output_MAC_86_27, I28=>output_MAC_86_28, I29=>output_MAC_86_29, I30=>output_MAC_86_30, I31=>output_MAC_86_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_86);

	mux_row_87: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_87_0, I1=>output_MAC_87_1, I2=>output_MAC_87_2, I3=>output_MAC_87_3, I4=>output_MAC_87_4, I5=>output_MAC_87_5, I6=>output_MAC_87_6, I7=>output_MAC_87_7, I8=>output_MAC_87_8, I9=>output_MAC_87_9, I10=>output_MAC_87_10, I11=>output_MAC_87_11, I12=>output_MAC_87_12, I13=>output_MAC_87_13, I14=>output_MAC_87_14, I15=>output_MAC_87_15, I16=>output_MAC_87_16, I17=>output_MAC_87_17, I18=>output_MAC_87_18, I19=>output_MAC_87_19, I20=>output_MAC_87_20, I21=>output_MAC_87_21, I22=>output_MAC_87_22, I23=>output_MAC_87_23, I24=>output_MAC_87_24, I25=>output_MAC_87_25, I26=>output_MAC_87_26, I27=>output_MAC_87_27, I28=>output_MAC_87_28, I29=>output_MAC_87_29, I30=>output_MAC_87_30, I31=>output_MAC_87_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_87);

	mux_row_88: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_88_0, I1=>output_MAC_88_1, I2=>output_MAC_88_2, I3=>output_MAC_88_3, I4=>output_MAC_88_4, I5=>output_MAC_88_5, I6=>output_MAC_88_6, I7=>output_MAC_88_7, I8=>output_MAC_88_8, I9=>output_MAC_88_9, I10=>output_MAC_88_10, I11=>output_MAC_88_11, I12=>output_MAC_88_12, I13=>output_MAC_88_13, I14=>output_MAC_88_14, I15=>output_MAC_88_15, I16=>output_MAC_88_16, I17=>output_MAC_88_17, I18=>output_MAC_88_18, I19=>output_MAC_88_19, I20=>output_MAC_88_20, I21=>output_MAC_88_21, I22=>output_MAC_88_22, I23=>output_MAC_88_23, I24=>output_MAC_88_24, I25=>output_MAC_88_25, I26=>output_MAC_88_26, I27=>output_MAC_88_27, I28=>output_MAC_88_28, I29=>output_MAC_88_29, I30=>output_MAC_88_30, I31=>output_MAC_88_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_88);

	mux_row_89: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_89_0, I1=>output_MAC_89_1, I2=>output_MAC_89_2, I3=>output_MAC_89_3, I4=>output_MAC_89_4, I5=>output_MAC_89_5, I6=>output_MAC_89_6, I7=>output_MAC_89_7, I8=>output_MAC_89_8, I9=>output_MAC_89_9, I10=>output_MAC_89_10, I11=>output_MAC_89_11, I12=>output_MAC_89_12, I13=>output_MAC_89_13, I14=>output_MAC_89_14, I15=>output_MAC_89_15, I16=>output_MAC_89_16, I17=>output_MAC_89_17, I18=>output_MAC_89_18, I19=>output_MAC_89_19, I20=>output_MAC_89_20, I21=>output_MAC_89_21, I22=>output_MAC_89_22, I23=>output_MAC_89_23, I24=>output_MAC_89_24, I25=>output_MAC_89_25, I26=>output_MAC_89_26, I27=>output_MAC_89_27, I28=>output_MAC_89_28, I29=>output_MAC_89_29, I30=>output_MAC_89_30, I31=>output_MAC_89_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_89);

	mux_row_90: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_90_0, I1=>output_MAC_90_1, I2=>output_MAC_90_2, I3=>output_MAC_90_3, I4=>output_MAC_90_4, I5=>output_MAC_90_5, I6=>output_MAC_90_6, I7=>output_MAC_90_7, I8=>output_MAC_90_8, I9=>output_MAC_90_9, I10=>output_MAC_90_10, I11=>output_MAC_90_11, I12=>output_MAC_90_12, I13=>output_MAC_90_13, I14=>output_MAC_90_14, I15=>output_MAC_90_15, I16=>output_MAC_90_16, I17=>output_MAC_90_17, I18=>output_MAC_90_18, I19=>output_MAC_90_19, I20=>output_MAC_90_20, I21=>output_MAC_90_21, I22=>output_MAC_90_22, I23=>output_MAC_90_23, I24=>output_MAC_90_24, I25=>output_MAC_90_25, I26=>output_MAC_90_26, I27=>output_MAC_90_27, I28=>output_MAC_90_28, I29=>output_MAC_90_29, I30=>output_MAC_90_30, I31=>output_MAC_90_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_90);

	mux_row_91: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_91_0, I1=>output_MAC_91_1, I2=>output_MAC_91_2, I3=>output_MAC_91_3, I4=>output_MAC_91_4, I5=>output_MAC_91_5, I6=>output_MAC_91_6, I7=>output_MAC_91_7, I8=>output_MAC_91_8, I9=>output_MAC_91_9, I10=>output_MAC_91_10, I11=>output_MAC_91_11, I12=>output_MAC_91_12, I13=>output_MAC_91_13, I14=>output_MAC_91_14, I15=>output_MAC_91_15, I16=>output_MAC_91_16, I17=>output_MAC_91_17, I18=>output_MAC_91_18, I19=>output_MAC_91_19, I20=>output_MAC_91_20, I21=>output_MAC_91_21, I22=>output_MAC_91_22, I23=>output_MAC_91_23, I24=>output_MAC_91_24, I25=>output_MAC_91_25, I26=>output_MAC_91_26, I27=>output_MAC_91_27, I28=>output_MAC_91_28, I29=>output_MAC_91_29, I30=>output_MAC_91_30, I31=>output_MAC_91_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_91);

	mux_row_92: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_92_0, I1=>output_MAC_92_1, I2=>output_MAC_92_2, I3=>output_MAC_92_3, I4=>output_MAC_92_4, I5=>output_MAC_92_5, I6=>output_MAC_92_6, I7=>output_MAC_92_7, I8=>output_MAC_92_8, I9=>output_MAC_92_9, I10=>output_MAC_92_10, I11=>output_MAC_92_11, I12=>output_MAC_92_12, I13=>output_MAC_92_13, I14=>output_MAC_92_14, I15=>output_MAC_92_15, I16=>output_MAC_92_16, I17=>output_MAC_92_17, I18=>output_MAC_92_18, I19=>output_MAC_92_19, I20=>output_MAC_92_20, I21=>output_MAC_92_21, I22=>output_MAC_92_22, I23=>output_MAC_92_23, I24=>output_MAC_92_24, I25=>output_MAC_92_25, I26=>output_MAC_92_26, I27=>output_MAC_92_27, I28=>output_MAC_92_28, I29=>output_MAC_92_29, I30=>output_MAC_92_30, I31=>output_MAC_92_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_92);

	mux_row_93: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_93_0, I1=>output_MAC_93_1, I2=>output_MAC_93_2, I3=>output_MAC_93_3, I4=>output_MAC_93_4, I5=>output_MAC_93_5, I6=>output_MAC_93_6, I7=>output_MAC_93_7, I8=>output_MAC_93_8, I9=>output_MAC_93_9, I10=>output_MAC_93_10, I11=>output_MAC_93_11, I12=>output_MAC_93_12, I13=>output_MAC_93_13, I14=>output_MAC_93_14, I15=>output_MAC_93_15, I16=>output_MAC_93_16, I17=>output_MAC_93_17, I18=>output_MAC_93_18, I19=>output_MAC_93_19, I20=>output_MAC_93_20, I21=>output_MAC_93_21, I22=>output_MAC_93_22, I23=>output_MAC_93_23, I24=>output_MAC_93_24, I25=>output_MAC_93_25, I26=>output_MAC_93_26, I27=>output_MAC_93_27, I28=>output_MAC_93_28, I29=>output_MAC_93_29, I30=>output_MAC_93_30, I31=>output_MAC_93_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_93);

	mux_row_94: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_94_0, I1=>output_MAC_94_1, I2=>output_MAC_94_2, I3=>output_MAC_94_3, I4=>output_MAC_94_4, I5=>output_MAC_94_5, I6=>output_MAC_94_6, I7=>output_MAC_94_7, I8=>output_MAC_94_8, I9=>output_MAC_94_9, I10=>output_MAC_94_10, I11=>output_MAC_94_11, I12=>output_MAC_94_12, I13=>output_MAC_94_13, I14=>output_MAC_94_14, I15=>output_MAC_94_15, I16=>output_MAC_94_16, I17=>output_MAC_94_17, I18=>output_MAC_94_18, I19=>output_MAC_94_19, I20=>output_MAC_94_20, I21=>output_MAC_94_21, I22=>output_MAC_94_22, I23=>output_MAC_94_23, I24=>output_MAC_94_24, I25=>output_MAC_94_25, I26=>output_MAC_94_26, I27=>output_MAC_94_27, I28=>output_MAC_94_28, I29=>output_MAC_94_29, I30=>output_MAC_94_30, I31=>output_MAC_94_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_94);

	mux_row_95: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_95_0, I1=>output_MAC_95_1, I2=>output_MAC_95_2, I3=>output_MAC_95_3, I4=>output_MAC_95_4, I5=>output_MAC_95_5, I6=>output_MAC_95_6, I7=>output_MAC_95_7, I8=>output_MAC_95_8, I9=>output_MAC_95_9, I10=>output_MAC_95_10, I11=>output_MAC_95_11, I12=>output_MAC_95_12, I13=>output_MAC_95_13, I14=>output_MAC_95_14, I15=>output_MAC_95_15, I16=>output_MAC_95_16, I17=>output_MAC_95_17, I18=>output_MAC_95_18, I19=>output_MAC_95_19, I20=>output_MAC_95_20, I21=>output_MAC_95_21, I22=>output_MAC_95_22, I23=>output_MAC_95_23, I24=>output_MAC_95_24, I25=>output_MAC_95_25, I26=>output_MAC_95_26, I27=>output_MAC_95_27, I28=>output_MAC_95_28, I29=>output_MAC_95_29, I30=>output_MAC_95_30, I31=>output_MAC_95_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_95);

	mux_row_96: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_96_0, I1=>output_MAC_96_1, I2=>output_MAC_96_2, I3=>output_MAC_96_3, I4=>output_MAC_96_4, I5=>output_MAC_96_5, I6=>output_MAC_96_6, I7=>output_MAC_96_7, I8=>output_MAC_96_8, I9=>output_MAC_96_9, I10=>output_MAC_96_10, I11=>output_MAC_96_11, I12=>output_MAC_96_12, I13=>output_MAC_96_13, I14=>output_MAC_96_14, I15=>output_MAC_96_15, I16=>output_MAC_96_16, I17=>output_MAC_96_17, I18=>output_MAC_96_18, I19=>output_MAC_96_19, I20=>output_MAC_96_20, I21=>output_MAC_96_21, I22=>output_MAC_96_22, I23=>output_MAC_96_23, I24=>output_MAC_96_24, I25=>output_MAC_96_25, I26=>output_MAC_96_26, I27=>output_MAC_96_27, I28=>output_MAC_96_28, I29=>output_MAC_96_29, I30=>output_MAC_96_30, I31=>output_MAC_96_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_96);

	mux_row_97: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_97_0, I1=>output_MAC_97_1, I2=>output_MAC_97_2, I3=>output_MAC_97_3, I4=>output_MAC_97_4, I5=>output_MAC_97_5, I6=>output_MAC_97_6, I7=>output_MAC_97_7, I8=>output_MAC_97_8, I9=>output_MAC_97_9, I10=>output_MAC_97_10, I11=>output_MAC_97_11, I12=>output_MAC_97_12, I13=>output_MAC_97_13, I14=>output_MAC_97_14, I15=>output_MAC_97_15, I16=>output_MAC_97_16, I17=>output_MAC_97_17, I18=>output_MAC_97_18, I19=>output_MAC_97_19, I20=>output_MAC_97_20, I21=>output_MAC_97_21, I22=>output_MAC_97_22, I23=>output_MAC_97_23, I24=>output_MAC_97_24, I25=>output_MAC_97_25, I26=>output_MAC_97_26, I27=>output_MAC_97_27, I28=>output_MAC_97_28, I29=>output_MAC_97_29, I30=>output_MAC_97_30, I31=>output_MAC_97_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_97);

	mux_row_98: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_98_0, I1=>output_MAC_98_1, I2=>output_MAC_98_2, I3=>output_MAC_98_3, I4=>output_MAC_98_4, I5=>output_MAC_98_5, I6=>output_MAC_98_6, I7=>output_MAC_98_7, I8=>output_MAC_98_8, I9=>output_MAC_98_9, I10=>output_MAC_98_10, I11=>output_MAC_98_11, I12=>output_MAC_98_12, I13=>output_MAC_98_13, I14=>output_MAC_98_14, I15=>output_MAC_98_15, I16=>output_MAC_98_16, I17=>output_MAC_98_17, I18=>output_MAC_98_18, I19=>output_MAC_98_19, I20=>output_MAC_98_20, I21=>output_MAC_98_21, I22=>output_MAC_98_22, I23=>output_MAC_98_23, I24=>output_MAC_98_24, I25=>output_MAC_98_25, I26=>output_MAC_98_26, I27=>output_MAC_98_27, I28=>output_MAC_98_28, I29=>output_MAC_98_29, I30=>output_MAC_98_30, I31=>output_MAC_98_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_98);

	mux_row_99: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_99_0, I1=>output_MAC_99_1, I2=>output_MAC_99_2, I3=>output_MAC_99_3, I4=>output_MAC_99_4, I5=>output_MAC_99_5, I6=>output_MAC_99_6, I7=>output_MAC_99_7, I8=>output_MAC_99_8, I9=>output_MAC_99_9, I10=>output_MAC_99_10, I11=>output_MAC_99_11, I12=>output_MAC_99_12, I13=>output_MAC_99_13, I14=>output_MAC_99_14, I15=>output_MAC_99_15, I16=>output_MAC_99_16, I17=>output_MAC_99_17, I18=>output_MAC_99_18, I19=>output_MAC_99_19, I20=>output_MAC_99_20, I21=>output_MAC_99_21, I22=>output_MAC_99_22, I23=>output_MAC_99_23, I24=>output_MAC_99_24, I25=>output_MAC_99_25, I26=>output_MAC_99_26, I27=>output_MAC_99_27, I28=>output_MAC_99_28, I29=>output_MAC_99_29, I30=>output_MAC_99_30, I31=>output_MAC_99_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_99);

	mux_row_100: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_100_0, I1=>output_MAC_100_1, I2=>output_MAC_100_2, I3=>output_MAC_100_3, I4=>output_MAC_100_4, I5=>output_MAC_100_5, I6=>output_MAC_100_6, I7=>output_MAC_100_7, I8=>output_MAC_100_8, I9=>output_MAC_100_9, I10=>output_MAC_100_10, I11=>output_MAC_100_11, I12=>output_MAC_100_12, I13=>output_MAC_100_13, I14=>output_MAC_100_14, I15=>output_MAC_100_15, I16=>output_MAC_100_16, I17=>output_MAC_100_17, I18=>output_MAC_100_18, I19=>output_MAC_100_19, I20=>output_MAC_100_20, I21=>output_MAC_100_21, I22=>output_MAC_100_22, I23=>output_MAC_100_23, I24=>output_MAC_100_24, I25=>output_MAC_100_25, I26=>output_MAC_100_26, I27=>output_MAC_100_27, I28=>output_MAC_100_28, I29=>output_MAC_100_29, I30=>output_MAC_100_30, I31=>output_MAC_100_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_100);

	mux_row_101: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_101_0, I1=>output_MAC_101_1, I2=>output_MAC_101_2, I3=>output_MAC_101_3, I4=>output_MAC_101_4, I5=>output_MAC_101_5, I6=>output_MAC_101_6, I7=>output_MAC_101_7, I8=>output_MAC_101_8, I9=>output_MAC_101_9, I10=>output_MAC_101_10, I11=>output_MAC_101_11, I12=>output_MAC_101_12, I13=>output_MAC_101_13, I14=>output_MAC_101_14, I15=>output_MAC_101_15, I16=>output_MAC_101_16, I17=>output_MAC_101_17, I18=>output_MAC_101_18, I19=>output_MAC_101_19, I20=>output_MAC_101_20, I21=>output_MAC_101_21, I22=>output_MAC_101_22, I23=>output_MAC_101_23, I24=>output_MAC_101_24, I25=>output_MAC_101_25, I26=>output_MAC_101_26, I27=>output_MAC_101_27, I28=>output_MAC_101_28, I29=>output_MAC_101_29, I30=>output_MAC_101_30, I31=>output_MAC_101_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_101);

	mux_row_102: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_102_0, I1=>output_MAC_102_1, I2=>output_MAC_102_2, I3=>output_MAC_102_3, I4=>output_MAC_102_4, I5=>output_MAC_102_5, I6=>output_MAC_102_6, I7=>output_MAC_102_7, I8=>output_MAC_102_8, I9=>output_MAC_102_9, I10=>output_MAC_102_10, I11=>output_MAC_102_11, I12=>output_MAC_102_12, I13=>output_MAC_102_13, I14=>output_MAC_102_14, I15=>output_MAC_102_15, I16=>output_MAC_102_16, I17=>output_MAC_102_17, I18=>output_MAC_102_18, I19=>output_MAC_102_19, I20=>output_MAC_102_20, I21=>output_MAC_102_21, I22=>output_MAC_102_22, I23=>output_MAC_102_23, I24=>output_MAC_102_24, I25=>output_MAC_102_25, I26=>output_MAC_102_26, I27=>output_MAC_102_27, I28=>output_MAC_102_28, I29=>output_MAC_102_29, I30=>output_MAC_102_30, I31=>output_MAC_102_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_102);

	mux_row_103: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_103_0, I1=>output_MAC_103_1, I2=>output_MAC_103_2, I3=>output_MAC_103_3, I4=>output_MAC_103_4, I5=>output_MAC_103_5, I6=>output_MAC_103_6, I7=>output_MAC_103_7, I8=>output_MAC_103_8, I9=>output_MAC_103_9, I10=>output_MAC_103_10, I11=>output_MAC_103_11, I12=>output_MAC_103_12, I13=>output_MAC_103_13, I14=>output_MAC_103_14, I15=>output_MAC_103_15, I16=>output_MAC_103_16, I17=>output_MAC_103_17, I18=>output_MAC_103_18, I19=>output_MAC_103_19, I20=>output_MAC_103_20, I21=>output_MAC_103_21, I22=>output_MAC_103_22, I23=>output_MAC_103_23, I24=>output_MAC_103_24, I25=>output_MAC_103_25, I26=>output_MAC_103_26, I27=>output_MAC_103_27, I28=>output_MAC_103_28, I29=>output_MAC_103_29, I30=>output_MAC_103_30, I31=>output_MAC_103_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_103);

	mux_row_104: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_104_0, I1=>output_MAC_104_1, I2=>output_MAC_104_2, I3=>output_MAC_104_3, I4=>output_MAC_104_4, I5=>output_MAC_104_5, I6=>output_MAC_104_6, I7=>output_MAC_104_7, I8=>output_MAC_104_8, I9=>output_MAC_104_9, I10=>output_MAC_104_10, I11=>output_MAC_104_11, I12=>output_MAC_104_12, I13=>output_MAC_104_13, I14=>output_MAC_104_14, I15=>output_MAC_104_15, I16=>output_MAC_104_16, I17=>output_MAC_104_17, I18=>output_MAC_104_18, I19=>output_MAC_104_19, I20=>output_MAC_104_20, I21=>output_MAC_104_21, I22=>output_MAC_104_22, I23=>output_MAC_104_23, I24=>output_MAC_104_24, I25=>output_MAC_104_25, I26=>output_MAC_104_26, I27=>output_MAC_104_27, I28=>output_MAC_104_28, I29=>output_MAC_104_29, I30=>output_MAC_104_30, I31=>output_MAC_104_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_104);

	mux_row_105: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_105_0, I1=>output_MAC_105_1, I2=>output_MAC_105_2, I3=>output_MAC_105_3, I4=>output_MAC_105_4, I5=>output_MAC_105_5, I6=>output_MAC_105_6, I7=>output_MAC_105_7, I8=>output_MAC_105_8, I9=>output_MAC_105_9, I10=>output_MAC_105_10, I11=>output_MAC_105_11, I12=>output_MAC_105_12, I13=>output_MAC_105_13, I14=>output_MAC_105_14, I15=>output_MAC_105_15, I16=>output_MAC_105_16, I17=>output_MAC_105_17, I18=>output_MAC_105_18, I19=>output_MAC_105_19, I20=>output_MAC_105_20, I21=>output_MAC_105_21, I22=>output_MAC_105_22, I23=>output_MAC_105_23, I24=>output_MAC_105_24, I25=>output_MAC_105_25, I26=>output_MAC_105_26, I27=>output_MAC_105_27, I28=>output_MAC_105_28, I29=>output_MAC_105_29, I30=>output_MAC_105_30, I31=>output_MAC_105_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_105);

	mux_row_106: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_106_0, I1=>output_MAC_106_1, I2=>output_MAC_106_2, I3=>output_MAC_106_3, I4=>output_MAC_106_4, I5=>output_MAC_106_5, I6=>output_MAC_106_6, I7=>output_MAC_106_7, I8=>output_MAC_106_8, I9=>output_MAC_106_9, I10=>output_MAC_106_10, I11=>output_MAC_106_11, I12=>output_MAC_106_12, I13=>output_MAC_106_13, I14=>output_MAC_106_14, I15=>output_MAC_106_15, I16=>output_MAC_106_16, I17=>output_MAC_106_17, I18=>output_MAC_106_18, I19=>output_MAC_106_19, I20=>output_MAC_106_20, I21=>output_MAC_106_21, I22=>output_MAC_106_22, I23=>output_MAC_106_23, I24=>output_MAC_106_24, I25=>output_MAC_106_25, I26=>output_MAC_106_26, I27=>output_MAC_106_27, I28=>output_MAC_106_28, I29=>output_MAC_106_29, I30=>output_MAC_106_30, I31=>output_MAC_106_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_106);

	mux_row_107: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_107_0, I1=>output_MAC_107_1, I2=>output_MAC_107_2, I3=>output_MAC_107_3, I4=>output_MAC_107_4, I5=>output_MAC_107_5, I6=>output_MAC_107_6, I7=>output_MAC_107_7, I8=>output_MAC_107_8, I9=>output_MAC_107_9, I10=>output_MAC_107_10, I11=>output_MAC_107_11, I12=>output_MAC_107_12, I13=>output_MAC_107_13, I14=>output_MAC_107_14, I15=>output_MAC_107_15, I16=>output_MAC_107_16, I17=>output_MAC_107_17, I18=>output_MAC_107_18, I19=>output_MAC_107_19, I20=>output_MAC_107_20, I21=>output_MAC_107_21, I22=>output_MAC_107_22, I23=>output_MAC_107_23, I24=>output_MAC_107_24, I25=>output_MAC_107_25, I26=>output_MAC_107_26, I27=>output_MAC_107_27, I28=>output_MAC_107_28, I29=>output_MAC_107_29, I30=>output_MAC_107_30, I31=>output_MAC_107_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_107);

	mux_row_108: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_108_0, I1=>output_MAC_108_1, I2=>output_MAC_108_2, I3=>output_MAC_108_3, I4=>output_MAC_108_4, I5=>output_MAC_108_5, I6=>output_MAC_108_6, I7=>output_MAC_108_7, I8=>output_MAC_108_8, I9=>output_MAC_108_9, I10=>output_MAC_108_10, I11=>output_MAC_108_11, I12=>output_MAC_108_12, I13=>output_MAC_108_13, I14=>output_MAC_108_14, I15=>output_MAC_108_15, I16=>output_MAC_108_16, I17=>output_MAC_108_17, I18=>output_MAC_108_18, I19=>output_MAC_108_19, I20=>output_MAC_108_20, I21=>output_MAC_108_21, I22=>output_MAC_108_22, I23=>output_MAC_108_23, I24=>output_MAC_108_24, I25=>output_MAC_108_25, I26=>output_MAC_108_26, I27=>output_MAC_108_27, I28=>output_MAC_108_28, I29=>output_MAC_108_29, I30=>output_MAC_108_30, I31=>output_MAC_108_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_108);

	mux_row_109: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_109_0, I1=>output_MAC_109_1, I2=>output_MAC_109_2, I3=>output_MAC_109_3, I4=>output_MAC_109_4, I5=>output_MAC_109_5, I6=>output_MAC_109_6, I7=>output_MAC_109_7, I8=>output_MAC_109_8, I9=>output_MAC_109_9, I10=>output_MAC_109_10, I11=>output_MAC_109_11, I12=>output_MAC_109_12, I13=>output_MAC_109_13, I14=>output_MAC_109_14, I15=>output_MAC_109_15, I16=>output_MAC_109_16, I17=>output_MAC_109_17, I18=>output_MAC_109_18, I19=>output_MAC_109_19, I20=>output_MAC_109_20, I21=>output_MAC_109_21, I22=>output_MAC_109_22, I23=>output_MAC_109_23, I24=>output_MAC_109_24, I25=>output_MAC_109_25, I26=>output_MAC_109_26, I27=>output_MAC_109_27, I28=>output_MAC_109_28, I29=>output_MAC_109_29, I30=>output_MAC_109_30, I31=>output_MAC_109_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_109);

	mux_row_110: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_110_0, I1=>output_MAC_110_1, I2=>output_MAC_110_2, I3=>output_MAC_110_3, I4=>output_MAC_110_4, I5=>output_MAC_110_5, I6=>output_MAC_110_6, I7=>output_MAC_110_7, I8=>output_MAC_110_8, I9=>output_MAC_110_9, I10=>output_MAC_110_10, I11=>output_MAC_110_11, I12=>output_MAC_110_12, I13=>output_MAC_110_13, I14=>output_MAC_110_14, I15=>output_MAC_110_15, I16=>output_MAC_110_16, I17=>output_MAC_110_17, I18=>output_MAC_110_18, I19=>output_MAC_110_19, I20=>output_MAC_110_20, I21=>output_MAC_110_21, I22=>output_MAC_110_22, I23=>output_MAC_110_23, I24=>output_MAC_110_24, I25=>output_MAC_110_25, I26=>output_MAC_110_26, I27=>output_MAC_110_27, I28=>output_MAC_110_28, I29=>output_MAC_110_29, I30=>output_MAC_110_30, I31=>output_MAC_110_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_110);

	mux_row_111: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_111_0, I1=>output_MAC_111_1, I2=>output_MAC_111_2, I3=>output_MAC_111_3, I4=>output_MAC_111_4, I5=>output_MAC_111_5, I6=>output_MAC_111_6, I7=>output_MAC_111_7, I8=>output_MAC_111_8, I9=>output_MAC_111_9, I10=>output_MAC_111_10, I11=>output_MAC_111_11, I12=>output_MAC_111_12, I13=>output_MAC_111_13, I14=>output_MAC_111_14, I15=>output_MAC_111_15, I16=>output_MAC_111_16, I17=>output_MAC_111_17, I18=>output_MAC_111_18, I19=>output_MAC_111_19, I20=>output_MAC_111_20, I21=>output_MAC_111_21, I22=>output_MAC_111_22, I23=>output_MAC_111_23, I24=>output_MAC_111_24, I25=>output_MAC_111_25, I26=>output_MAC_111_26, I27=>output_MAC_111_27, I28=>output_MAC_111_28, I29=>output_MAC_111_29, I30=>output_MAC_111_30, I31=>output_MAC_111_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_111);

	mux_row_112: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_112_0, I1=>output_MAC_112_1, I2=>output_MAC_112_2, I3=>output_MAC_112_3, I4=>output_MAC_112_4, I5=>output_MAC_112_5, I6=>output_MAC_112_6, I7=>output_MAC_112_7, I8=>output_MAC_112_8, I9=>output_MAC_112_9, I10=>output_MAC_112_10, I11=>output_MAC_112_11, I12=>output_MAC_112_12, I13=>output_MAC_112_13, I14=>output_MAC_112_14, I15=>output_MAC_112_15, I16=>output_MAC_112_16, I17=>output_MAC_112_17, I18=>output_MAC_112_18, I19=>output_MAC_112_19, I20=>output_MAC_112_20, I21=>output_MAC_112_21, I22=>output_MAC_112_22, I23=>output_MAC_112_23, I24=>output_MAC_112_24, I25=>output_MAC_112_25, I26=>output_MAC_112_26, I27=>output_MAC_112_27, I28=>output_MAC_112_28, I29=>output_MAC_112_29, I30=>output_MAC_112_30, I31=>output_MAC_112_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_112);

	mux_row_113: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_113_0, I1=>output_MAC_113_1, I2=>output_MAC_113_2, I3=>output_MAC_113_3, I4=>output_MAC_113_4, I5=>output_MAC_113_5, I6=>output_MAC_113_6, I7=>output_MAC_113_7, I8=>output_MAC_113_8, I9=>output_MAC_113_9, I10=>output_MAC_113_10, I11=>output_MAC_113_11, I12=>output_MAC_113_12, I13=>output_MAC_113_13, I14=>output_MAC_113_14, I15=>output_MAC_113_15, I16=>output_MAC_113_16, I17=>output_MAC_113_17, I18=>output_MAC_113_18, I19=>output_MAC_113_19, I20=>output_MAC_113_20, I21=>output_MAC_113_21, I22=>output_MAC_113_22, I23=>output_MAC_113_23, I24=>output_MAC_113_24, I25=>output_MAC_113_25, I26=>output_MAC_113_26, I27=>output_MAC_113_27, I28=>output_MAC_113_28, I29=>output_MAC_113_29, I30=>output_MAC_113_30, I31=>output_MAC_113_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_113);

	mux_row_114: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_114_0, I1=>output_MAC_114_1, I2=>output_MAC_114_2, I3=>output_MAC_114_3, I4=>output_MAC_114_4, I5=>output_MAC_114_5, I6=>output_MAC_114_6, I7=>output_MAC_114_7, I8=>output_MAC_114_8, I9=>output_MAC_114_9, I10=>output_MAC_114_10, I11=>output_MAC_114_11, I12=>output_MAC_114_12, I13=>output_MAC_114_13, I14=>output_MAC_114_14, I15=>output_MAC_114_15, I16=>output_MAC_114_16, I17=>output_MAC_114_17, I18=>output_MAC_114_18, I19=>output_MAC_114_19, I20=>output_MAC_114_20, I21=>output_MAC_114_21, I22=>output_MAC_114_22, I23=>output_MAC_114_23, I24=>output_MAC_114_24, I25=>output_MAC_114_25, I26=>output_MAC_114_26, I27=>output_MAC_114_27, I28=>output_MAC_114_28, I29=>output_MAC_114_29, I30=>output_MAC_114_30, I31=>output_MAC_114_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_114);

	mux_row_115: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_115_0, I1=>output_MAC_115_1, I2=>output_MAC_115_2, I3=>output_MAC_115_3, I4=>output_MAC_115_4, I5=>output_MAC_115_5, I6=>output_MAC_115_6, I7=>output_MAC_115_7, I8=>output_MAC_115_8, I9=>output_MAC_115_9, I10=>output_MAC_115_10, I11=>output_MAC_115_11, I12=>output_MAC_115_12, I13=>output_MAC_115_13, I14=>output_MAC_115_14, I15=>output_MAC_115_15, I16=>output_MAC_115_16, I17=>output_MAC_115_17, I18=>output_MAC_115_18, I19=>output_MAC_115_19, I20=>output_MAC_115_20, I21=>output_MAC_115_21, I22=>output_MAC_115_22, I23=>output_MAC_115_23, I24=>output_MAC_115_24, I25=>output_MAC_115_25, I26=>output_MAC_115_26, I27=>output_MAC_115_27, I28=>output_MAC_115_28, I29=>output_MAC_115_29, I30=>output_MAC_115_30, I31=>output_MAC_115_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_115);

	mux_row_116: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_116_0, I1=>output_MAC_116_1, I2=>output_MAC_116_2, I3=>output_MAC_116_3, I4=>output_MAC_116_4, I5=>output_MAC_116_5, I6=>output_MAC_116_6, I7=>output_MAC_116_7, I8=>output_MAC_116_8, I9=>output_MAC_116_9, I10=>output_MAC_116_10, I11=>output_MAC_116_11, I12=>output_MAC_116_12, I13=>output_MAC_116_13, I14=>output_MAC_116_14, I15=>output_MAC_116_15, I16=>output_MAC_116_16, I17=>output_MAC_116_17, I18=>output_MAC_116_18, I19=>output_MAC_116_19, I20=>output_MAC_116_20, I21=>output_MAC_116_21, I22=>output_MAC_116_22, I23=>output_MAC_116_23, I24=>output_MAC_116_24, I25=>output_MAC_116_25, I26=>output_MAC_116_26, I27=>output_MAC_116_27, I28=>output_MAC_116_28, I29=>output_MAC_116_29, I30=>output_MAC_116_30, I31=>output_MAC_116_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_116);

	mux_row_117: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_117_0, I1=>output_MAC_117_1, I2=>output_MAC_117_2, I3=>output_MAC_117_3, I4=>output_MAC_117_4, I5=>output_MAC_117_5, I6=>output_MAC_117_6, I7=>output_MAC_117_7, I8=>output_MAC_117_8, I9=>output_MAC_117_9, I10=>output_MAC_117_10, I11=>output_MAC_117_11, I12=>output_MAC_117_12, I13=>output_MAC_117_13, I14=>output_MAC_117_14, I15=>output_MAC_117_15, I16=>output_MAC_117_16, I17=>output_MAC_117_17, I18=>output_MAC_117_18, I19=>output_MAC_117_19, I20=>output_MAC_117_20, I21=>output_MAC_117_21, I22=>output_MAC_117_22, I23=>output_MAC_117_23, I24=>output_MAC_117_24, I25=>output_MAC_117_25, I26=>output_MAC_117_26, I27=>output_MAC_117_27, I28=>output_MAC_117_28, I29=>output_MAC_117_29, I30=>output_MAC_117_30, I31=>output_MAC_117_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_117);

	mux_row_118: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_118_0, I1=>output_MAC_118_1, I2=>output_MAC_118_2, I3=>output_MAC_118_3, I4=>output_MAC_118_4, I5=>output_MAC_118_5, I6=>output_MAC_118_6, I7=>output_MAC_118_7, I8=>output_MAC_118_8, I9=>output_MAC_118_9, I10=>output_MAC_118_10, I11=>output_MAC_118_11, I12=>output_MAC_118_12, I13=>output_MAC_118_13, I14=>output_MAC_118_14, I15=>output_MAC_118_15, I16=>output_MAC_118_16, I17=>output_MAC_118_17, I18=>output_MAC_118_18, I19=>output_MAC_118_19, I20=>output_MAC_118_20, I21=>output_MAC_118_21, I22=>output_MAC_118_22, I23=>output_MAC_118_23, I24=>output_MAC_118_24, I25=>output_MAC_118_25, I26=>output_MAC_118_26, I27=>output_MAC_118_27, I28=>output_MAC_118_28, I29=>output_MAC_118_29, I30=>output_MAC_118_30, I31=>output_MAC_118_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_118);

	mux_row_119: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_119_0, I1=>output_MAC_119_1, I2=>output_MAC_119_2, I3=>output_MAC_119_3, I4=>output_MAC_119_4, I5=>output_MAC_119_5, I6=>output_MAC_119_6, I7=>output_MAC_119_7, I8=>output_MAC_119_8, I9=>output_MAC_119_9, I10=>output_MAC_119_10, I11=>output_MAC_119_11, I12=>output_MAC_119_12, I13=>output_MAC_119_13, I14=>output_MAC_119_14, I15=>output_MAC_119_15, I16=>output_MAC_119_16, I17=>output_MAC_119_17, I18=>output_MAC_119_18, I19=>output_MAC_119_19, I20=>output_MAC_119_20, I21=>output_MAC_119_21, I22=>output_MAC_119_22, I23=>output_MAC_119_23, I24=>output_MAC_119_24, I25=>output_MAC_119_25, I26=>output_MAC_119_26, I27=>output_MAC_119_27, I28=>output_MAC_119_28, I29=>output_MAC_119_29, I30=>output_MAC_119_30, I31=>output_MAC_119_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_119);

	mux_row_120: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_120_0, I1=>output_MAC_120_1, I2=>output_MAC_120_2, I3=>output_MAC_120_3, I4=>output_MAC_120_4, I5=>output_MAC_120_5, I6=>output_MAC_120_6, I7=>output_MAC_120_7, I8=>output_MAC_120_8, I9=>output_MAC_120_9, I10=>output_MAC_120_10, I11=>output_MAC_120_11, I12=>output_MAC_120_12, I13=>output_MAC_120_13, I14=>output_MAC_120_14, I15=>output_MAC_120_15, I16=>output_MAC_120_16, I17=>output_MAC_120_17, I18=>output_MAC_120_18, I19=>output_MAC_120_19, I20=>output_MAC_120_20, I21=>output_MAC_120_21, I22=>output_MAC_120_22, I23=>output_MAC_120_23, I24=>output_MAC_120_24, I25=>output_MAC_120_25, I26=>output_MAC_120_26, I27=>output_MAC_120_27, I28=>output_MAC_120_28, I29=>output_MAC_120_29, I30=>output_MAC_120_30, I31=>output_MAC_120_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_120);

	mux_row_121: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_121_0, I1=>output_MAC_121_1, I2=>output_MAC_121_2, I3=>output_MAC_121_3, I4=>output_MAC_121_4, I5=>output_MAC_121_5, I6=>output_MAC_121_6, I7=>output_MAC_121_7, I8=>output_MAC_121_8, I9=>output_MAC_121_9, I10=>output_MAC_121_10, I11=>output_MAC_121_11, I12=>output_MAC_121_12, I13=>output_MAC_121_13, I14=>output_MAC_121_14, I15=>output_MAC_121_15, I16=>output_MAC_121_16, I17=>output_MAC_121_17, I18=>output_MAC_121_18, I19=>output_MAC_121_19, I20=>output_MAC_121_20, I21=>output_MAC_121_21, I22=>output_MAC_121_22, I23=>output_MAC_121_23, I24=>output_MAC_121_24, I25=>output_MAC_121_25, I26=>output_MAC_121_26, I27=>output_MAC_121_27, I28=>output_MAC_121_28, I29=>output_MAC_121_29, I30=>output_MAC_121_30, I31=>output_MAC_121_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_121);

	mux_row_122: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_122_0, I1=>output_MAC_122_1, I2=>output_MAC_122_2, I3=>output_MAC_122_3, I4=>output_MAC_122_4, I5=>output_MAC_122_5, I6=>output_MAC_122_6, I7=>output_MAC_122_7, I8=>output_MAC_122_8, I9=>output_MAC_122_9, I10=>output_MAC_122_10, I11=>output_MAC_122_11, I12=>output_MAC_122_12, I13=>output_MAC_122_13, I14=>output_MAC_122_14, I15=>output_MAC_122_15, I16=>output_MAC_122_16, I17=>output_MAC_122_17, I18=>output_MAC_122_18, I19=>output_MAC_122_19, I20=>output_MAC_122_20, I21=>output_MAC_122_21, I22=>output_MAC_122_22, I23=>output_MAC_122_23, I24=>output_MAC_122_24, I25=>output_MAC_122_25, I26=>output_MAC_122_26, I27=>output_MAC_122_27, I28=>output_MAC_122_28, I29=>output_MAC_122_29, I30=>output_MAC_122_30, I31=>output_MAC_122_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_122);

	mux_row_123: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_123_0, I1=>output_MAC_123_1, I2=>output_MAC_123_2, I3=>output_MAC_123_3, I4=>output_MAC_123_4, I5=>output_MAC_123_5, I6=>output_MAC_123_6, I7=>output_MAC_123_7, I8=>output_MAC_123_8, I9=>output_MAC_123_9, I10=>output_MAC_123_10, I11=>output_MAC_123_11, I12=>output_MAC_123_12, I13=>output_MAC_123_13, I14=>output_MAC_123_14, I15=>output_MAC_123_15, I16=>output_MAC_123_16, I17=>output_MAC_123_17, I18=>output_MAC_123_18, I19=>output_MAC_123_19, I20=>output_MAC_123_20, I21=>output_MAC_123_21, I22=>output_MAC_123_22, I23=>output_MAC_123_23, I24=>output_MAC_123_24, I25=>output_MAC_123_25, I26=>output_MAC_123_26, I27=>output_MAC_123_27, I28=>output_MAC_123_28, I29=>output_MAC_123_29, I30=>output_MAC_123_30, I31=>output_MAC_123_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_123);

	mux_row_124: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_124_0, I1=>output_MAC_124_1, I2=>output_MAC_124_2, I3=>output_MAC_124_3, I4=>output_MAC_124_4, I5=>output_MAC_124_5, I6=>output_MAC_124_6, I7=>output_MAC_124_7, I8=>output_MAC_124_8, I9=>output_MAC_124_9, I10=>output_MAC_124_10, I11=>output_MAC_124_11, I12=>output_MAC_124_12, I13=>output_MAC_124_13, I14=>output_MAC_124_14, I15=>output_MAC_124_15, I16=>output_MAC_124_16, I17=>output_MAC_124_17, I18=>output_MAC_124_18, I19=>output_MAC_124_19, I20=>output_MAC_124_20, I21=>output_MAC_124_21, I22=>output_MAC_124_22, I23=>output_MAC_124_23, I24=>output_MAC_124_24, I25=>output_MAC_124_25, I26=>output_MAC_124_26, I27=>output_MAC_124_27, I28=>output_MAC_124_28, I29=>output_MAC_124_29, I30=>output_MAC_124_30, I31=>output_MAC_124_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_124);

	mux_row_125: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_125_0, I1=>output_MAC_125_1, I2=>output_MAC_125_2, I3=>output_MAC_125_3, I4=>output_MAC_125_4, I5=>output_MAC_125_5, I6=>output_MAC_125_6, I7=>output_MAC_125_7, I8=>output_MAC_125_8, I9=>output_MAC_125_9, I10=>output_MAC_125_10, I11=>output_MAC_125_11, I12=>output_MAC_125_12, I13=>output_MAC_125_13, I14=>output_MAC_125_14, I15=>output_MAC_125_15, I16=>output_MAC_125_16, I17=>output_MAC_125_17, I18=>output_MAC_125_18, I19=>output_MAC_125_19, I20=>output_MAC_125_20, I21=>output_MAC_125_21, I22=>output_MAC_125_22, I23=>output_MAC_125_23, I24=>output_MAC_125_24, I25=>output_MAC_125_25, I26=>output_MAC_125_26, I27=>output_MAC_125_27, I28=>output_MAC_125_28, I29=>output_MAC_125_29, I30=>output_MAC_125_30, I31=>output_MAC_125_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_125);

	mux_row_126: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_126_0, I1=>output_MAC_126_1, I2=>output_MAC_126_2, I3=>output_MAC_126_3, I4=>output_MAC_126_4, I5=>output_MAC_126_5, I6=>output_MAC_126_6, I7=>output_MAC_126_7, I8=>output_MAC_126_8, I9=>output_MAC_126_9, I10=>output_MAC_126_10, I11=>output_MAC_126_11, I12=>output_MAC_126_12, I13=>output_MAC_126_13, I14=>output_MAC_126_14, I15=>output_MAC_126_15, I16=>output_MAC_126_16, I17=>output_MAC_126_17, I18=>output_MAC_126_18, I19=>output_MAC_126_19, I20=>output_MAC_126_20, I21=>output_MAC_126_21, I22=>output_MAC_126_22, I23=>output_MAC_126_23, I24=>output_MAC_126_24, I25=>output_MAC_126_25, I26=>output_MAC_126_26, I27=>output_MAC_126_27, I28=>output_MAC_126_28, I29=>output_MAC_126_29, I30=>output_MAC_126_30, I31=>output_MAC_126_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_126);

	mux_row_127: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_127_0, I1=>output_MAC_127_1, I2=>output_MAC_127_2, I3=>output_MAC_127_3, I4=>output_MAC_127_4, I5=>output_MAC_127_5, I6=>output_MAC_127_6, I7=>output_MAC_127_7, I8=>output_MAC_127_8, I9=>output_MAC_127_9, I10=>output_MAC_127_10, I11=>output_MAC_127_11, I12=>output_MAC_127_12, I13=>output_MAC_127_13, I14=>output_MAC_127_14, I15=>output_MAC_127_15, I16=>output_MAC_127_16, I17=>output_MAC_127_17, I18=>output_MAC_127_18, I19=>output_MAC_127_19, I20=>output_MAC_127_20, I21=>output_MAC_127_21, I22=>output_MAC_127_22, I23=>output_MAC_127_23, I24=>output_MAC_127_24, I25=>output_MAC_127_25, I26=>output_MAC_127_26, I27=>output_MAC_127_27, I28=>output_MAC_127_28, I29=>output_MAC_127_29, I30=>output_MAC_127_30, I31=>output_MAC_127_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_127);

	output_row_0_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_0, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_0);
	output_row_1_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_1, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_1);
	output_row_2_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_2, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_2);
	output_row_3_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_3, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_3);
	output_row_4_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_4, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_4);
	output_row_5_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_5, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_5);
	output_row_6_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_6, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_6);
	output_row_7_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_7, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_7);
	output_row_8_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_8, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_8);
	output_row_9_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_9, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_9);
	output_row_10_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_10, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_10);
	output_row_11_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_11, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_11);
	output_row_12_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_12, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_12);
	output_row_13_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_13, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_13);
	output_row_14_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_14, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_14);
	output_row_15_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_15, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_15);
	output_row_16_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_16, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_16);
	output_row_17_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_17, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_17);
	output_row_18_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_18, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_18);
	output_row_19_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_19, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_19);
	output_row_20_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_20, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_20);
	output_row_21_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_21, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_21);
	output_row_22_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_22, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_22);
	output_row_23_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_23, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_23);
	output_row_24_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_24, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_24);
	output_row_25_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_25, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_25);
	output_row_26_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_26, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_26);
	output_row_27_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_27, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_27);
	output_row_28_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_28, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_28);
	output_row_29_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_29, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_29);
	output_row_30_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_30, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_30);
	output_row_31_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_31, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_31);
	output_row_32_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_32, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_32);
	output_row_33_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_33, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_33);
	output_row_34_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_34, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_34);
	output_row_35_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_35, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_35);
	output_row_36_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_36, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_36);
	output_row_37_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_37, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_37);
	output_row_38_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_38, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_38);
	output_row_39_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_39, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_39);
	output_row_40_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_40, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_40);
	output_row_41_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_41, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_41);
	output_row_42_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_42, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_42);
	output_row_43_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_43, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_43);
	output_row_44_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_44, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_44);
	output_row_45_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_45, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_45);
	output_row_46_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_46, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_46);
	output_row_47_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_47, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_47);
	output_row_48_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_48, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_48);
	output_row_49_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_49, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_49);
	output_row_50_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_50, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_50);
	output_row_51_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_51, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_51);
	output_row_52_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_52, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_52);
	output_row_53_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_53, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_53);
	output_row_54_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_54, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_54);
	output_row_55_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_55, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_55);
	output_row_56_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_56, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_56);
	output_row_57_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_57, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_57);
	output_row_58_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_58, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_58);
	output_row_59_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_59, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_59);
	output_row_60_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_60, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_60);
	output_row_61_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_61, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_61);
	output_row_62_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_62, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_62);
	output_row_63_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_63, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_63);
	output_row_64_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_64, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_64);
	output_row_65_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_65, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_65);
	output_row_66_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_66, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_66);
	output_row_67_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_67, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_67);
	output_row_68_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_68, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_68);
	output_row_69_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_69, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_69);
	output_row_70_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_70, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_70);
	output_row_71_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_71, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_71);
	output_row_72_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_72, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_72);
	output_row_73_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_73, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_73);
	output_row_74_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_74, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_74);
	output_row_75_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_75, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_75);
	output_row_76_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_76, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_76);
	output_row_77_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_77, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_77);
	output_row_78_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_78, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_78);
	output_row_79_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_79, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_79);
	output_row_80_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_80, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_80);
	output_row_81_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_81, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_81);
	output_row_82_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_82, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_82);
	output_row_83_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_83, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_83);
	output_row_84_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_84, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_84);
	output_row_85_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_85, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_85);
	output_row_86_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_86, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_86);
	output_row_87_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_87, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_87);
	output_row_88_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_88, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_88);
	output_row_89_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_89, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_89);
	output_row_90_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_90, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_90);
	output_row_91_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_91, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_91);
	output_row_92_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_92, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_92);
	output_row_93_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_93, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_93);
	output_row_94_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_94, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_94);
	output_row_95_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_95, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_95);
	output_row_96_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_96, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_96);
	output_row_97_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_97, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_97);
	output_row_98_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_98, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_98);
	output_row_99_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_99, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_99);
	output_row_100_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_100, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_100);
	output_row_101_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_101, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_101);
	output_row_102_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_102, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_102);
	output_row_103_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_103, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_103);
	output_row_104_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_104, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_104);
	output_row_105_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_105, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_105);
	output_row_106_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_106, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_106);
	output_row_107_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_107, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_107);
	output_row_108_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_108, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_108);
	output_row_109_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_109, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_109);
	output_row_110_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_110, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_110);
	output_row_111_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_111, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_111);
	output_row_112_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_112, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_112);
	output_row_113_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_113, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_113);
	output_row_114_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_114, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_114);
	output_row_115_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_115, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_115);
	output_row_116_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_116, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_116);
	output_row_117_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_117, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_117);
	output_row_118_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_118, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_118);
	output_row_119_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_119, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_119);
	output_row_120_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_120, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_120);
	output_row_121_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_121, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_121);
	output_row_122_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_122, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_122);
	output_row_123_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_123, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_123);
	output_row_124_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_124, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_124);
	output_row_125_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_125, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_125);
	output_row_126_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_126, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_126);
	output_row_127_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_127, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_127);

END behaviour;
