
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mux_768to1_nbit IS
GENERIC(
	N : POSITIVE := 2
);
PORT (I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, 
	I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, 
	I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, 
	I30, I31, I32, I33, I34, I35, I36, I37, I38, I39, 
	I40, I41, I42, I43, I44, I45, I46, I47, I48, I49, 
	I50, I51, I52, I53, I54, I55, I56, I57, I58, I59, 
	I60, I61, I62, I63, I64, I65, I66, I67, I68, I69, 
	I70, I71, I72, I73, I74, I75, I76, I77, I78, I79, 
	I80, I81, I82, I83, I84, I85, I86, I87, I88, I89, 
	I90, I91, I92, I93, I94, I95, I96, I97, I98, I99, 
	I100, I101, I102, I103, I104, I105, I106, I107, I108, I109, 
	I110, I111, I112, I113, I114, I115, I116, I117, I118, I119, 
	I120, I121, I122, I123, I124, I125, I126, I127, I128, I129, 
	I130, I131, I132, I133, I134, I135, I136, I137, I138, I139, 
	I140, I141, I142, I143, I144, I145, I146, I147, I148, I149, 
	I150, I151, I152, I153, I154, I155, I156, I157, I158, I159, 
	I160, I161, I162, I163, I164, I165, I166, I167, I168, I169, 
	I170, I171, I172, I173, I174, I175, I176, I177, I178, I179, 
	I180, I181, I182, I183, I184, I185, I186, I187, I188, I189, 
	I190, I191, I192, I193, I194, I195, I196, I197, I198, I199, 
	I200, I201, I202, I203, I204, I205, I206, I207, I208, I209, 
	I210, I211, I212, I213, I214, I215, I216, I217, I218, I219, 
	I220, I221, I222, I223, I224, I225, I226, I227, I228, I229, 
	I230, I231, I232, I233, I234, I235, I236, I237, I238, I239, 
	I240, I241, I242, I243, I244, I245, I246, I247, I248, I249, 
	I250, I251, I252, I253, I254, I255, I256, I257, I258, I259, 
	I260, I261, I262, I263, I264, I265, I266, I267, I268, I269, 
	I270, I271, I272, I273, I274, I275, I276, I277, I278, I279, 
	I280, I281, I282, I283, I284, I285, I286, I287, I288, I289, 
	I290, I291, I292, I293, I294, I295, I296, I297, I298, I299, 
	I300, I301, I302, I303, I304, I305, I306, I307, I308, I309, 
	I310, I311, I312, I313, I314, I315, I316, I317, I318, I319, 
	I320, I321, I322, I323, I324, I325, I326, I327, I328, I329, 
	I330, I331, I332, I333, I334, I335, I336, I337, I338, I339, 
	I340, I341, I342, I343, I344, I345, I346, I347, I348, I349, 
	I350, I351, I352, I353, I354, I355, I356, I357, I358, I359, 
	I360, I361, I362, I363, I364, I365, I366, I367, I368, I369, 
	I370, I371, I372, I373, I374, I375, I376, I377, I378, I379, 
	I380, I381, I382, I383, I384, I385, I386, I387, I388, I389, 
	I390, I391, I392, I393, I394, I395, I396, I397, I398, I399, 
	I400, I401, I402, I403, I404, I405, I406, I407, I408, I409, 
	I410, I411, I412, I413, I414, I415, I416, I417, I418, I419, 
	I420, I421, I422, I423, I424, I425, I426, I427, I428, I429, 
	I430, I431, I432, I433, I434, I435, I436, I437, I438, I439, 
	I440, I441, I442, I443, I444, I445, I446, I447, I448, I449, 
	I450, I451, I452, I453, I454, I455, I456, I457, I458, I459, 
	I460, I461, I462, I463, I464, I465, I466, I467, I468, I469, 
	I470, I471, I472, I473, I474, I475, I476, I477, I478, I479, 
	I480, I481, I482, I483, I484, I485, I486, I487, I488, I489, 
	I490, I491, I492, I493, I494, I495, I496, I497, I498, I499, 
	I500, I501, I502, I503, I504, I505, I506, I507, I508, I509, 
	I510, I511, I512, I513, I514, I515, I516, I517, I518, I519, 
	I520, I521, I522, I523, I524, I525, I526, I527, I528, I529, 
	I530, I531, I532, I533, I534, I535, I536, I537, I538, I539, 
	I540, I541, I542, I543, I544, I545, I546, I547, I548, I549, 
	I550, I551, I552, I553, I554, I555, I556, I557, I558, I559, 
	I560, I561, I562, I563, I564, I565, I566, I567, I568, I569, 
	I570, I571, I572, I573, I574, I575, I576, I577, I578, I579, 
	I580, I581, I582, I583, I584, I585, I586, I587, I588, I589, 
	I590, I591, I592, I593, I594, I595, I596, I597, I598, I599, 
	I600, I601, I602, I603, I604, I605, I606, I607, I608, I609, 
	I610, I611, I612, I613, I614, I615, I616, I617, I618, I619, 
	I620, I621, I622, I623, I624, I625, I626, I627, I628, I629, 
	I630, I631, I632, I633, I634, I635, I636, I637, I638, I639, 
	I640, I641, I642, I643, I644, I645, I646, I647, I648, I649, 
	I650, I651, I652, I653, I654, I655, I656, I657, I658, I659, 
	I660, I661, I662, I663, I664, I665, I666, I667, I668, I669, 
	I670, I671, I672, I673, I674, I675, I676, I677, I678, I679, 
	I680, I681, I682, I683, I684, I685, I686, I687, I688, I689, 
	I690, I691, I692, I693, I694, I695, I696, I697, I698, I699, 
	I700, I701, I702, I703, I704, I705, I706, I707, I708, I709, 
	I710, I711, I712, I713, I714, I715, I716, I717, I718, I719, 
	I720, I721, I722, I723, I724, I725, I726, I727, I728, I729, 
	I730, I731, I732, I733, I734, I735, I736, I737, I738, I739, 
	I740, I741, I742, I743, I744, I745, I746, I747, I748, I749, 
	I750, I751, I752, I753, I754, I755, I756, I757, I758, I759, 
	I760, I761, I762, I763, I764, I765, I766, I767: IN STD_LOGIC_VECTOR(N-1 downto 0);
	SEL_mux: IN STD_LOGIC_VECTOR(9 downto 0);
	O: OUT STD_LOGIC_VECTOR(N-1 downto 0)
);
END mux_768to1_nbit;

ARCHITECTURE behaviour OF  mux_768to1_nbit IS

COMPONENT mux_4to1_nbit_base IS
	GENERIC ( N : POSITIVE :=1);
	PORT( I0, I1, I2, I3: IN STD_LOGIC_VECTOR(N-1 downto 0);
		SEL  : IN STD_LOGIC_VECTOR(1 downto 0);
		O    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
END COMPONENT;

COMPONENT mux_2to1_nbit_base IS
GENERIC ( N : POSITIVE :=1
);
PORT( 
	I0, I1: IN STD_LOGIC_VECTOR(N-1 downto 0);
	SEL  : IN STD_LOGIC;
	O    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
		 );
END COMPONENT;


SIGNAL output_mux_0_0: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_1: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_2: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_3: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_4: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_5: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_6: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_7: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_8: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_9: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_10: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_11: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_12: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_13: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_14: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_15: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_16: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_17: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_18: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_19: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_20: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_21: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_22: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_23: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_24: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_25: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_26: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_27: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_28: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_29: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_30: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_31: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_32: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_33: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_34: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_35: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_36: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_37: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_38: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_39: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_40: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_41: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_42: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_43: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_44: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_45: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_46: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_47: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_48: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_49: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_50: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_51: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_52: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_53: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_54: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_55: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_56: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_57: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_58: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_59: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_60: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_61: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_62: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_63: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_64: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_65: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_66: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_67: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_68: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_69: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_70: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_71: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_72: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_73: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_74: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_75: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_76: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_77: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_78: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_79: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_80: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_81: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_82: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_83: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_84: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_85: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_86: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_87: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_88: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_89: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_90: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_91: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_92: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_93: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_94: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_95: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_96: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_97: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_98: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_99: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_100: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_101: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_102: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_103: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_104: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_105: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_106: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_107: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_108: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_109: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_110: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_111: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_112: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_113: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_114: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_115: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_116: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_117: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_118: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_119: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_120: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_121: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_122: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_123: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_124: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_125: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_126: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_127: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_128: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_129: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_130: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_131: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_132: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_133: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_134: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_135: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_136: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_137: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_138: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_139: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_140: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_141: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_142: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_143: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_144: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_145: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_146: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_147: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_148: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_149: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_150: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_151: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_152: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_153: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_154: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_155: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_156: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_157: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_158: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_159: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_160: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_161: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_162: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_163: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_164: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_165: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_166: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_167: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_168: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_169: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_170: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_171: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_172: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_173: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_174: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_175: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_176: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_177: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_178: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_179: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_180: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_181: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_182: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_183: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_184: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_185: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_186: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_187: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_188: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_189: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_190: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_0_191: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_0: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_1: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_2: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_3: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_4: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_5: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_6: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_7: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_8: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_9: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_10: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_11: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_12: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_13: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_14: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_15: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_16: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_17: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_18: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_19: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_20: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_21: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_22: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_23: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_24: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_25: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_26: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_27: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_28: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_29: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_30: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_31: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_32: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_33: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_34: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_35: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_36: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_37: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_38: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_39: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_40: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_41: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_42: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_43: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_44: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_45: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_46: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_1_47: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_0: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_1: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_2: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_3: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_4: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_5: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_6: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_7: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_8: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_9: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_10: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_2_11: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_3_0: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_3_1: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_3_2: STD_LOGIC_VECTOR(N-1 downto 0);
SIGNAL output_mux_4_0: STD_LOGIC_VECTOR(N-1 downto 0);

BEGIN

mux_0_0: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I0, I1=>I1, I2=>I2, I3=>I3, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_0);
mux_0_1: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I4, I1=>I5, I2=>I6, I3=>I7, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_1);
mux_0_2: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I8, I1=>I9, I2=>I10, I3=>I11, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_2);
mux_0_3: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I12, I1=>I13, I2=>I14, I3=>I15, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_3);
mux_0_4: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I16, I1=>I17, I2=>I18, I3=>I19, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_4);
mux_0_5: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I20, I1=>I21, I2=>I22, I3=>I23, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_5);
mux_0_6: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I24, I1=>I25, I2=>I26, I3=>I27, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_6);
mux_0_7: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I28, I1=>I29, I2=>I30, I3=>I31, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_7);
mux_0_8: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I32, I1=>I33, I2=>I34, I3=>I35, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_8);
mux_0_9: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I36, I1=>I37, I2=>I38, I3=>I39, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_9);
mux_0_10: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I40, I1=>I41, I2=>I42, I3=>I43, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_10);
mux_0_11: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I44, I1=>I45, I2=>I46, I3=>I47, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_11);
mux_0_12: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I48, I1=>I49, I2=>I50, I3=>I51, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_12);
mux_0_13: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I52, I1=>I53, I2=>I54, I3=>I55, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_13);
mux_0_14: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I56, I1=>I57, I2=>I58, I3=>I59, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_14);
mux_0_15: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I60, I1=>I61, I2=>I62, I3=>I63, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_15);
mux_0_16: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I64, I1=>I65, I2=>I66, I3=>I67, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_16);
mux_0_17: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I68, I1=>I69, I2=>I70, I3=>I71, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_17);
mux_0_18: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I72, I1=>I73, I2=>I74, I3=>I75, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_18);
mux_0_19: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I76, I1=>I77, I2=>I78, I3=>I79, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_19);
mux_0_20: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I80, I1=>I81, I2=>I82, I3=>I83, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_20);
mux_0_21: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I84, I1=>I85, I2=>I86, I3=>I87, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_21);
mux_0_22: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I88, I1=>I89, I2=>I90, I3=>I91, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_22);
mux_0_23: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I92, I1=>I93, I2=>I94, I3=>I95, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_23);
mux_0_24: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I96, I1=>I97, I2=>I98, I3=>I99, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_24);
mux_0_25: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I100, I1=>I101, I2=>I102, I3=>I103, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_25);
mux_0_26: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I104, I1=>I105, I2=>I106, I3=>I107, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_26);
mux_0_27: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I108, I1=>I109, I2=>I110, I3=>I111, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_27);
mux_0_28: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I112, I1=>I113, I2=>I114, I3=>I115, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_28);
mux_0_29: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I116, I1=>I117, I2=>I118, I3=>I119, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_29);
mux_0_30: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I120, I1=>I121, I2=>I122, I3=>I123, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_30);
mux_0_31: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I124, I1=>I125, I2=>I126, I3=>I127, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_31);
mux_0_32: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I128, I1=>I129, I2=>I130, I3=>I131, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_32);
mux_0_33: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I132, I1=>I133, I2=>I134, I3=>I135, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_33);
mux_0_34: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I136, I1=>I137, I2=>I138, I3=>I139, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_34);
mux_0_35: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I140, I1=>I141, I2=>I142, I3=>I143, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_35);
mux_0_36: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I144, I1=>I145, I2=>I146, I3=>I147, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_36);
mux_0_37: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I148, I1=>I149, I2=>I150, I3=>I151, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_37);
mux_0_38: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I152, I1=>I153, I2=>I154, I3=>I155, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_38);
mux_0_39: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I156, I1=>I157, I2=>I158, I3=>I159, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_39);
mux_0_40: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I160, I1=>I161, I2=>I162, I3=>I163, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_40);
mux_0_41: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I164, I1=>I165, I2=>I166, I3=>I167, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_41);
mux_0_42: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I168, I1=>I169, I2=>I170, I3=>I171, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_42);
mux_0_43: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I172, I1=>I173, I2=>I174, I3=>I175, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_43);
mux_0_44: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I176, I1=>I177, I2=>I178, I3=>I179, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_44);
mux_0_45: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I180, I1=>I181, I2=>I182, I3=>I183, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_45);
mux_0_46: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I184, I1=>I185, I2=>I186, I3=>I187, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_46);
mux_0_47: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I188, I1=>I189, I2=>I190, I3=>I191, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_47);
mux_0_48: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I192, I1=>I193, I2=>I194, I3=>I195, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_48);
mux_0_49: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I196, I1=>I197, I2=>I198, I3=>I199, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_49);
mux_0_50: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I200, I1=>I201, I2=>I202, I3=>I203, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_50);
mux_0_51: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I204, I1=>I205, I2=>I206, I3=>I207, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_51);
mux_0_52: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I208, I1=>I209, I2=>I210, I3=>I211, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_52);
mux_0_53: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I212, I1=>I213, I2=>I214, I3=>I215, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_53);
mux_0_54: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I216, I1=>I217, I2=>I218, I3=>I219, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_54);
mux_0_55: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I220, I1=>I221, I2=>I222, I3=>I223, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_55);
mux_0_56: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I224, I1=>I225, I2=>I226, I3=>I227, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_56);
mux_0_57: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I228, I1=>I229, I2=>I230, I3=>I231, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_57);
mux_0_58: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I232, I1=>I233, I2=>I234, I3=>I235, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_58);
mux_0_59: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I236, I1=>I237, I2=>I238, I3=>I239, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_59);
mux_0_60: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I240, I1=>I241, I2=>I242, I3=>I243, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_60);
mux_0_61: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I244, I1=>I245, I2=>I246, I3=>I247, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_61);
mux_0_62: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I248, I1=>I249, I2=>I250, I3=>I251, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_62);
mux_0_63: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I252, I1=>I253, I2=>I254, I3=>I255, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_63);
mux_0_64: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I256, I1=>I257, I2=>I258, I3=>I259, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_64);
mux_0_65: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I260, I1=>I261, I2=>I262, I3=>I263, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_65);
mux_0_66: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I264, I1=>I265, I2=>I266, I3=>I267, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_66);
mux_0_67: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I268, I1=>I269, I2=>I270, I3=>I271, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_67);
mux_0_68: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I272, I1=>I273, I2=>I274, I3=>I275, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_68);
mux_0_69: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I276, I1=>I277, I2=>I278, I3=>I279, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_69);
mux_0_70: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I280, I1=>I281, I2=>I282, I3=>I283, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_70);
mux_0_71: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I284, I1=>I285, I2=>I286, I3=>I287, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_71);
mux_0_72: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I288, I1=>I289, I2=>I290, I3=>I291, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_72);
mux_0_73: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I292, I1=>I293, I2=>I294, I3=>I295, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_73);
mux_0_74: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I296, I1=>I297, I2=>I298, I3=>I299, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_74);
mux_0_75: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I300, I1=>I301, I2=>I302, I3=>I303, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_75);
mux_0_76: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I304, I1=>I305, I2=>I306, I3=>I307, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_76);
mux_0_77: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I308, I1=>I309, I2=>I310, I3=>I311, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_77);
mux_0_78: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I312, I1=>I313, I2=>I314, I3=>I315, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_78);
mux_0_79: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I316, I1=>I317, I2=>I318, I3=>I319, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_79);
mux_0_80: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I320, I1=>I321, I2=>I322, I3=>I323, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_80);
mux_0_81: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I324, I1=>I325, I2=>I326, I3=>I327, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_81);
mux_0_82: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I328, I1=>I329, I2=>I330, I3=>I331, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_82);
mux_0_83: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I332, I1=>I333, I2=>I334, I3=>I335, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_83);
mux_0_84: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I336, I1=>I337, I2=>I338, I3=>I339, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_84);
mux_0_85: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I340, I1=>I341, I2=>I342, I3=>I343, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_85);
mux_0_86: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I344, I1=>I345, I2=>I346, I3=>I347, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_86);
mux_0_87: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I348, I1=>I349, I2=>I350, I3=>I351, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_87);
mux_0_88: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I352, I1=>I353, I2=>I354, I3=>I355, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_88);
mux_0_89: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I356, I1=>I357, I2=>I358, I3=>I359, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_89);
mux_0_90: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I360, I1=>I361, I2=>I362, I3=>I363, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_90);
mux_0_91: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I364, I1=>I365, I2=>I366, I3=>I367, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_91);
mux_0_92: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I368, I1=>I369, I2=>I370, I3=>I371, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_92);
mux_0_93: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I372, I1=>I373, I2=>I374, I3=>I375, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_93);
mux_0_94: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I376, I1=>I377, I2=>I378, I3=>I379, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_94);
mux_0_95: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I380, I1=>I381, I2=>I382, I3=>I383, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_95);
mux_0_96: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I384, I1=>I385, I2=>I386, I3=>I387, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_96);
mux_0_97: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I388, I1=>I389, I2=>I390, I3=>I391, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_97);
mux_0_98: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I392, I1=>I393, I2=>I394, I3=>I395, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_98);
mux_0_99: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I396, I1=>I397, I2=>I398, I3=>I399, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_99);
mux_0_100: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I400, I1=>I401, I2=>I402, I3=>I403, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_100);
mux_0_101: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I404, I1=>I405, I2=>I406, I3=>I407, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_101);
mux_0_102: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I408, I1=>I409, I2=>I410, I3=>I411, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_102);
mux_0_103: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I412, I1=>I413, I2=>I414, I3=>I415, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_103);
mux_0_104: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I416, I1=>I417, I2=>I418, I3=>I419, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_104);
mux_0_105: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I420, I1=>I421, I2=>I422, I3=>I423, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_105);
mux_0_106: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I424, I1=>I425, I2=>I426, I3=>I427, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_106);
mux_0_107: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I428, I1=>I429, I2=>I430, I3=>I431, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_107);
mux_0_108: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I432, I1=>I433, I2=>I434, I3=>I435, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_108);
mux_0_109: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I436, I1=>I437, I2=>I438, I3=>I439, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_109);
mux_0_110: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I440, I1=>I441, I2=>I442, I3=>I443, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_110);
mux_0_111: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I444, I1=>I445, I2=>I446, I3=>I447, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_111);
mux_0_112: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I448, I1=>I449, I2=>I450, I3=>I451, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_112);
mux_0_113: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I452, I1=>I453, I2=>I454, I3=>I455, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_113);
mux_0_114: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I456, I1=>I457, I2=>I458, I3=>I459, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_114);
mux_0_115: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I460, I1=>I461, I2=>I462, I3=>I463, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_115);
mux_0_116: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I464, I1=>I465, I2=>I466, I3=>I467, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_116);
mux_0_117: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I468, I1=>I469, I2=>I470, I3=>I471, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_117);
mux_0_118: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I472, I1=>I473, I2=>I474, I3=>I475, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_118);
mux_0_119: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I476, I1=>I477, I2=>I478, I3=>I479, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_119);
mux_0_120: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I480, I1=>I481, I2=>I482, I3=>I483, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_120);
mux_0_121: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I484, I1=>I485, I2=>I486, I3=>I487, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_121);
mux_0_122: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I488, I1=>I489, I2=>I490, I3=>I491, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_122);
mux_0_123: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I492, I1=>I493, I2=>I494, I3=>I495, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_123);
mux_0_124: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I496, I1=>I497, I2=>I498, I3=>I499, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_124);
mux_0_125: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I500, I1=>I501, I2=>I502, I3=>I503, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_125);
mux_0_126: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I504, I1=>I505, I2=>I506, I3=>I507, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_126);
mux_0_127: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I508, I1=>I509, I2=>I510, I3=>I511, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_127);
mux_0_128: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I512, I1=>I513, I2=>I514, I3=>I515, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_128);
mux_0_129: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I516, I1=>I517, I2=>I518, I3=>I519, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_129);
mux_0_130: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I520, I1=>I521, I2=>I522, I3=>I523, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_130);
mux_0_131: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I524, I1=>I525, I2=>I526, I3=>I527, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_131);
mux_0_132: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I528, I1=>I529, I2=>I530, I3=>I531, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_132);
mux_0_133: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I532, I1=>I533, I2=>I534, I3=>I535, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_133);
mux_0_134: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I536, I1=>I537, I2=>I538, I3=>I539, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_134);
mux_0_135: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I540, I1=>I541, I2=>I542, I3=>I543, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_135);
mux_0_136: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I544, I1=>I545, I2=>I546, I3=>I547, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_136);
mux_0_137: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I548, I1=>I549, I2=>I550, I3=>I551, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_137);
mux_0_138: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I552, I1=>I553, I2=>I554, I3=>I555, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_138);
mux_0_139: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I556, I1=>I557, I2=>I558, I3=>I559, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_139);
mux_0_140: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I560, I1=>I561, I2=>I562, I3=>I563, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_140);
mux_0_141: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I564, I1=>I565, I2=>I566, I3=>I567, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_141);
mux_0_142: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I568, I1=>I569, I2=>I570, I3=>I571, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_142);
mux_0_143: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I572, I1=>I573, I2=>I574, I3=>I575, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_143);
mux_0_144: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I576, I1=>I577, I2=>I578, I3=>I579, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_144);
mux_0_145: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I580, I1=>I581, I2=>I582, I3=>I583, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_145);
mux_0_146: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I584, I1=>I585, I2=>I586, I3=>I587, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_146);
mux_0_147: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I588, I1=>I589, I2=>I590, I3=>I591, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_147);
mux_0_148: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I592, I1=>I593, I2=>I594, I3=>I595, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_148);
mux_0_149: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I596, I1=>I597, I2=>I598, I3=>I599, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_149);
mux_0_150: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I600, I1=>I601, I2=>I602, I3=>I603, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_150);
mux_0_151: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I604, I1=>I605, I2=>I606, I3=>I607, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_151);
mux_0_152: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I608, I1=>I609, I2=>I610, I3=>I611, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_152);
mux_0_153: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I612, I1=>I613, I2=>I614, I3=>I615, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_153);
mux_0_154: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I616, I1=>I617, I2=>I618, I3=>I619, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_154);
mux_0_155: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I620, I1=>I621, I2=>I622, I3=>I623, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_155);
mux_0_156: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I624, I1=>I625, I2=>I626, I3=>I627, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_156);
mux_0_157: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I628, I1=>I629, I2=>I630, I3=>I631, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_157);
mux_0_158: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I632, I1=>I633, I2=>I634, I3=>I635, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_158);
mux_0_159: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I636, I1=>I637, I2=>I638, I3=>I639, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_159);
mux_0_160: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I640, I1=>I641, I2=>I642, I3=>I643, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_160);
mux_0_161: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I644, I1=>I645, I2=>I646, I3=>I647, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_161);
mux_0_162: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I648, I1=>I649, I2=>I650, I3=>I651, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_162);
mux_0_163: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I652, I1=>I653, I2=>I654, I3=>I655, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_163);
mux_0_164: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I656, I1=>I657, I2=>I658, I3=>I659, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_164);
mux_0_165: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I660, I1=>I661, I2=>I662, I3=>I663, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_165);
mux_0_166: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I664, I1=>I665, I2=>I666, I3=>I667, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_166);
mux_0_167: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I668, I1=>I669, I2=>I670, I3=>I671, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_167);
mux_0_168: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I672, I1=>I673, I2=>I674, I3=>I675, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_168);
mux_0_169: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I676, I1=>I677, I2=>I678, I3=>I679, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_169);
mux_0_170: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I680, I1=>I681, I2=>I682, I3=>I683, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_170);
mux_0_171: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I684, I1=>I685, I2=>I686, I3=>I687, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_171);
mux_0_172: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I688, I1=>I689, I2=>I690, I3=>I691, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_172);
mux_0_173: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I692, I1=>I693, I2=>I694, I3=>I695, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_173);
mux_0_174: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I696, I1=>I697, I2=>I698, I3=>I699, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_174);
mux_0_175: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I700, I1=>I701, I2=>I702, I3=>I703, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_175);
mux_0_176: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I704, I1=>I705, I2=>I706, I3=>I707, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_176);
mux_0_177: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I708, I1=>I709, I2=>I710, I3=>I711, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_177);
mux_0_178: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I712, I1=>I713, I2=>I714, I3=>I715, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_178);
mux_0_179: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I716, I1=>I717, I2=>I718, I3=>I719, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_179);
mux_0_180: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I720, I1=>I721, I2=>I722, I3=>I723, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_180);
mux_0_181: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I724, I1=>I725, I2=>I726, I3=>I727, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_181);
mux_0_182: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I728, I1=>I729, I2=>I730, I3=>I731, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_182);
mux_0_183: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I732, I1=>I733, I2=>I734, I3=>I735, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_183);
mux_0_184: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I736, I1=>I737, I2=>I738, I3=>I739, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_184);
mux_0_185: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I740, I1=>I741, I2=>I742, I3=>I743, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_185);
mux_0_186: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I744, I1=>I745, I2=>I746, I3=>I747, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_186);
mux_0_187: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I748, I1=>I749, I2=>I750, I3=>I751, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_187);
mux_0_188: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I752, I1=>I753, I2=>I754, I3=>I755, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_188);
mux_0_189: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I756, I1=>I757, I2=>I758, I3=>I759, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_189);
mux_0_190: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I760, I1=>I761, I2=>I762, I3=>I763, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_190);
mux_0_191: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>I764, I1=>I765, I2=>I766, I3=>I767, SEL=>SEL_mux(1 downto 0), O=>output_mux_0_191);
mux_1_0: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_0, I1=>output_mux_0_1, I2=>output_mux_0_2, I3=>output_mux_0_3, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_0);
mux_1_1: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_4, I1=>output_mux_0_5, I2=>output_mux_0_6, I3=>output_mux_0_7, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_1);
mux_1_2: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_8, I1=>output_mux_0_9, I2=>output_mux_0_10, I3=>output_mux_0_11, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_2);
mux_1_3: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_12, I1=>output_mux_0_13, I2=>output_mux_0_14, I3=>output_mux_0_15, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_3);
mux_1_4: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_16, I1=>output_mux_0_17, I2=>output_mux_0_18, I3=>output_mux_0_19, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_4);
mux_1_5: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_20, I1=>output_mux_0_21, I2=>output_mux_0_22, I3=>output_mux_0_23, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_5);
mux_1_6: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_24, I1=>output_mux_0_25, I2=>output_mux_0_26, I3=>output_mux_0_27, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_6);
mux_1_7: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_28, I1=>output_mux_0_29, I2=>output_mux_0_30, I3=>output_mux_0_31, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_7);
mux_1_8: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_32, I1=>output_mux_0_33, I2=>output_mux_0_34, I3=>output_mux_0_35, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_8);
mux_1_9: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_36, I1=>output_mux_0_37, I2=>output_mux_0_38, I3=>output_mux_0_39, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_9);
mux_1_10: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_40, I1=>output_mux_0_41, I2=>output_mux_0_42, I3=>output_mux_0_43, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_10);
mux_1_11: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_44, I1=>output_mux_0_45, I2=>output_mux_0_46, I3=>output_mux_0_47, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_11);
mux_1_12: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_48, I1=>output_mux_0_49, I2=>output_mux_0_50, I3=>output_mux_0_51, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_12);
mux_1_13: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_52, I1=>output_mux_0_53, I2=>output_mux_0_54, I3=>output_mux_0_55, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_13);
mux_1_14: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_56, I1=>output_mux_0_57, I2=>output_mux_0_58, I3=>output_mux_0_59, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_14);
mux_1_15: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_60, I1=>output_mux_0_61, I2=>output_mux_0_62, I3=>output_mux_0_63, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_15);
mux_1_16: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_64, I1=>output_mux_0_65, I2=>output_mux_0_66, I3=>output_mux_0_67, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_16);
mux_1_17: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_68, I1=>output_mux_0_69, I2=>output_mux_0_70, I3=>output_mux_0_71, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_17);
mux_1_18: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_72, I1=>output_mux_0_73, I2=>output_mux_0_74, I3=>output_mux_0_75, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_18);
mux_1_19: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_76, I1=>output_mux_0_77, I2=>output_mux_0_78, I3=>output_mux_0_79, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_19);
mux_1_20: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_80, I1=>output_mux_0_81, I2=>output_mux_0_82, I3=>output_mux_0_83, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_20);
mux_1_21: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_84, I1=>output_mux_0_85, I2=>output_mux_0_86, I3=>output_mux_0_87, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_21);
mux_1_22: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_88, I1=>output_mux_0_89, I2=>output_mux_0_90, I3=>output_mux_0_91, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_22);
mux_1_23: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_92, I1=>output_mux_0_93, I2=>output_mux_0_94, I3=>output_mux_0_95, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_23);
mux_1_24: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_96, I1=>output_mux_0_97, I2=>output_mux_0_98, I3=>output_mux_0_99, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_24);
mux_1_25: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_100, I1=>output_mux_0_101, I2=>output_mux_0_102, I3=>output_mux_0_103, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_25);
mux_1_26: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_104, I1=>output_mux_0_105, I2=>output_mux_0_106, I3=>output_mux_0_107, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_26);
mux_1_27: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_108, I1=>output_mux_0_109, I2=>output_mux_0_110, I3=>output_mux_0_111, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_27);
mux_1_28: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_112, I1=>output_mux_0_113, I2=>output_mux_0_114, I3=>output_mux_0_115, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_28);
mux_1_29: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_116, I1=>output_mux_0_117, I2=>output_mux_0_118, I3=>output_mux_0_119, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_29);
mux_1_30: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_120, I1=>output_mux_0_121, I2=>output_mux_0_122, I3=>output_mux_0_123, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_30);
mux_1_31: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_124, I1=>output_mux_0_125, I2=>output_mux_0_126, I3=>output_mux_0_127, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_31);
mux_1_32: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_128, I1=>output_mux_0_129, I2=>output_mux_0_130, I3=>output_mux_0_131, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_32);
mux_1_33: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_132, I1=>output_mux_0_133, I2=>output_mux_0_134, I3=>output_mux_0_135, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_33);
mux_1_34: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_136, I1=>output_mux_0_137, I2=>output_mux_0_138, I3=>output_mux_0_139, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_34);
mux_1_35: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_140, I1=>output_mux_0_141, I2=>output_mux_0_142, I3=>output_mux_0_143, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_35);
mux_1_36: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_144, I1=>output_mux_0_145, I2=>output_mux_0_146, I3=>output_mux_0_147, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_36);
mux_1_37: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_148, I1=>output_mux_0_149, I2=>output_mux_0_150, I3=>output_mux_0_151, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_37);
mux_1_38: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_152, I1=>output_mux_0_153, I2=>output_mux_0_154, I3=>output_mux_0_155, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_38);
mux_1_39: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_156, I1=>output_mux_0_157, I2=>output_mux_0_158, I3=>output_mux_0_159, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_39);
mux_1_40: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_160, I1=>output_mux_0_161, I2=>output_mux_0_162, I3=>output_mux_0_163, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_40);
mux_1_41: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_164, I1=>output_mux_0_165, I2=>output_mux_0_166, I3=>output_mux_0_167, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_41);
mux_1_42: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_168, I1=>output_mux_0_169, I2=>output_mux_0_170, I3=>output_mux_0_171, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_42);
mux_1_43: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_172, I1=>output_mux_0_173, I2=>output_mux_0_174, I3=>output_mux_0_175, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_43);
mux_1_44: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_176, I1=>output_mux_0_177, I2=>output_mux_0_178, I3=>output_mux_0_179, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_44);
mux_1_45: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_180, I1=>output_mux_0_181, I2=>output_mux_0_182, I3=>output_mux_0_183, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_45);
mux_1_46: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_184, I1=>output_mux_0_185, I2=>output_mux_0_186, I3=>output_mux_0_187, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_46);
mux_1_47: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_0_188, I1=>output_mux_0_189, I2=>output_mux_0_190, I3=>output_mux_0_191, SEL=>SEL_mux(3 downto 2), O=>output_mux_1_47);
mux_2_0: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_0, I1=>output_mux_1_1, I2=>output_mux_1_2, I3=>output_mux_1_3, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_0);
mux_2_1: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_4, I1=>output_mux_1_5, I2=>output_mux_1_6, I3=>output_mux_1_7, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_1);
mux_2_2: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_8, I1=>output_mux_1_9, I2=>output_mux_1_10, I3=>output_mux_1_11, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_2);
mux_2_3: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_12, I1=>output_mux_1_13, I2=>output_mux_1_14, I3=>output_mux_1_15, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_3);
mux_2_4: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_16, I1=>output_mux_1_17, I2=>output_mux_1_18, I3=>output_mux_1_19, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_4);
mux_2_5: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_20, I1=>output_mux_1_21, I2=>output_mux_1_22, I3=>output_mux_1_23, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_5);
mux_2_6: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_24, I1=>output_mux_1_25, I2=>output_mux_1_26, I3=>output_mux_1_27, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_6);
mux_2_7: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_28, I1=>output_mux_1_29, I2=>output_mux_1_30, I3=>output_mux_1_31, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_7);
mux_2_8: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_32, I1=>output_mux_1_33, I2=>output_mux_1_34, I3=>output_mux_1_35, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_8);
mux_2_9: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_36, I1=>output_mux_1_37, I2=>output_mux_1_38, I3=>output_mux_1_39, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_9);
mux_2_10: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_40, I1=>output_mux_1_41, I2=>output_mux_1_42, I3=>output_mux_1_43, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_10);
mux_2_11: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_1_44, I1=>output_mux_1_45, I2=>output_mux_1_46, I3=>output_mux_1_47, SEL=>SEL_mux(5 downto 4), O=>output_mux_2_11);
mux_3_0: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_2_0, I1=>output_mux_2_1, I2=>output_mux_2_2, I3=>output_mux_2_3, SEL=>SEL_mux(7 downto 6), O=>output_mux_3_0);
mux_3_1: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_2_4, I1=>output_mux_2_5, I2=>output_mux_2_6, I3=>output_mux_2_7, SEL=>SEL_mux(7 downto 6), O=>output_mux_3_1);
mux_3_2: mux_4to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_2_8, I1=>output_mux_2_9, I2=>output_mux_2_10, I3=>output_mux_2_11, SEL=>SEL_mux(7 downto 6), O=>output_mux_3_2);

mux_4_0: mux_2to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_3_0, I1=>output_mux_3_1, SEL=>SEL_mux(8), O=>output_mux_4_0);

mux_5_0: mux_2to1_nbit_base GENERIC MAP(N=>N) PORT MAP(I0=>output_mux_4_0, I1=>output_mux_3_2, SEL=>SEL_mux(9), O=>O);

END behaviour;
