
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MAC_32x32_8_reg IS
PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7, input_row_8, input_row_9, 
	input_row_10, input_row_11, input_row_12, input_row_13, input_row_14, input_row_15, input_row_16, input_row_17, input_row_18, input_row_19, 
	input_row_20, input_row_21, input_row_22, input_row_23, input_row_24, input_row_25, input_row_26, input_row_27, input_row_28, input_row_29, 
	input_row_30, input_row_31: IN STD_LOGIC_VECTOR(7 downto 0);
	input_col_0, input_col_1, input_col_2, input_col_3, input_col_4, input_col_5, input_col_6, input_col_7, input_col_8, input_col_9, 
	input_col_10, input_col_11, input_col_12, input_col_13, input_col_14, input_col_15, input_col_16, input_col_17, input_col_18, input_col_19, 
	input_col_20, input_col_21, input_col_22, input_col_23, input_col_24, input_col_25, input_col_26, input_col_27, input_col_28, input_col_29, 
	input_col_30, input_col_31: IN STD_LOGIC_VECTOR(7 downto 0);
	SEL_mux: IN STD_LOGIC_VECTOR(4 downto 0);
	CLK, RST_n, ENABLE : IN STD_LOGIC;
	output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7, output_row_8, output_row_9, 
	output_row_10, output_row_11, output_row_12, output_row_13, output_row_14, output_row_15, output_row_16, output_row_17, output_row_18, output_row_19, 
	output_row_20, output_row_21, output_row_22, output_row_23, output_row_24, output_row_25, output_row_26, output_row_27, output_row_28, output_row_29, 
	output_row_30, output_row_31: OUT STD_LOGIC_VECTOR(31 downto 0)
);
END MAC_32x32_8_reg;

ARCHITECTURE behaviour OF  MAC_32x32_8_reg IS

	COMPONENT MAC IS
	GENERIC (data_size : POSITIVE := 2; 
	acc_size: POSITIVE := 16	);
	PORT( data_in_A, data_in_B  : IN STD_LOGIC_VECTOR(data_size-1 downto 0);
		CLK, RST_n, ENABLE 	: IN STD_LOGIC;
		data_out    			: OUT STD_LOGIC_VECTOR(acc_size-1 downto 0));
	END COMPONENT;

	COMPONENT mux_32to1_nbit IS
	GENERIC ( N : POSITIVE :=2);
	PORT(
		I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, 
		I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, 
		I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, 
		I30, I31: IN STD_LOGIC_VECTOR(N-1 downto 0);
		SEL_mux  : IN STD_LOGIC_VECTOR(4 downto 0);
		O    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
	END COMPONENT;

	COMPONENT regnbit IS
	GENERIC ( N : POSITIVE := 2);
	PORT(
		D    : IN STD_LOGIC_VECTOR(N-1 downto 0);
		CLK, RST_n, ENABLE : IN STD_LOGIC;
		Q    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
	END COMPONENT;

	COMPONENT ff IS
	PORT(
		D    : IN STD_LOGIC;
		CLK, RST_n, ENABLE : IN STD_LOGIC;
		Q    : OUT STD_LOGIC
	);
	END COMPONENT;

	SIGNAL reg_input_row_0, reg_input_row_1, reg_input_row_2, reg_input_row_3, reg_input_row_4, reg_input_row_5, reg_input_row_6, reg_input_row_7, reg_input_row_8, reg_input_row_9, 
		reg_input_row_10, reg_input_row_11, reg_input_row_12, reg_input_row_13, reg_input_row_14, reg_input_row_15, reg_input_row_16, reg_input_row_17, reg_input_row_18, reg_input_row_19, 
		reg_input_row_20, reg_input_row_21, reg_input_row_22, reg_input_row_23, reg_input_row_24, reg_input_row_25, reg_input_row_26, reg_input_row_27, reg_input_row_28, reg_input_row_29, 
		reg_input_row_30, reg_input_row_31: STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL reg_input_col_0, reg_input_col_1, reg_input_col_2, reg_input_col_3, reg_input_col_4, reg_input_col_5, reg_input_col_6, reg_input_col_7, reg_input_col_8, reg_input_col_9, 
		reg_input_col_10, reg_input_col_11, reg_input_col_12, reg_input_col_13, reg_input_col_14, reg_input_col_15, reg_input_col_16, reg_input_col_17, reg_input_col_18, reg_input_col_19, 
		reg_input_col_20, reg_input_col_21, reg_input_col_22, reg_input_col_23, reg_input_col_24, reg_input_col_25, reg_input_col_26, reg_input_col_27, reg_input_col_28, reg_input_col_29, 
		reg_input_col_30, reg_input_col_31: STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL reg_SEL_mux: STD_LOGIC_VECTOR(4 downto 0);
	SIGNAL reg_ENABLE_in, reg_ENABLE_out : STD_LOGIC;
	SIGNAL reg_output_row_0, reg_output_row_1, reg_output_row_2, reg_output_row_3, reg_output_row_4, reg_output_row_5, reg_output_row_6, reg_output_row_7, reg_output_row_8, reg_output_row_9, 
		reg_output_row_10, reg_output_row_11, reg_output_row_12, reg_output_row_13, reg_output_row_14, reg_output_row_15, reg_output_row_16, reg_output_row_17, reg_output_row_18, reg_output_row_19, 
		reg_output_row_20, reg_output_row_21, reg_output_row_22, reg_output_row_23, reg_output_row_24, reg_output_row_25, reg_output_row_26, reg_output_row_27, reg_output_row_28, reg_output_row_29, 
		reg_output_row_30, reg_output_row_31: STD_LOGIC_VECTOR(31 downto 0);

	SIGNAL output_MAC_0_0, output_MAC_0_1, output_MAC_0_2, output_MAC_0_3, output_MAC_0_4, output_MAC_0_5, output_MAC_0_6, output_MAC_0_7, output_MAC_0_8, output_MAC_0_9, 
		output_MAC_0_10, output_MAC_0_11, output_MAC_0_12, output_MAC_0_13, output_MAC_0_14, output_MAC_0_15, output_MAC_0_16, output_MAC_0_17, output_MAC_0_18, output_MAC_0_19, 
		output_MAC_0_20, output_MAC_0_21, output_MAC_0_22, output_MAC_0_23, output_MAC_0_24, output_MAC_0_25, output_MAC_0_26, output_MAC_0_27, output_MAC_0_28, output_MAC_0_29, 
		output_MAC_0_30, output_MAC_0_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_1_0, output_MAC_1_1, output_MAC_1_2, output_MAC_1_3, output_MAC_1_4, output_MAC_1_5, output_MAC_1_6, output_MAC_1_7, output_MAC_1_8, output_MAC_1_9, 
		output_MAC_1_10, output_MAC_1_11, output_MAC_1_12, output_MAC_1_13, output_MAC_1_14, output_MAC_1_15, output_MAC_1_16, output_MAC_1_17, output_MAC_1_18, output_MAC_1_19, 
		output_MAC_1_20, output_MAC_1_21, output_MAC_1_22, output_MAC_1_23, output_MAC_1_24, output_MAC_1_25, output_MAC_1_26, output_MAC_1_27, output_MAC_1_28, output_MAC_1_29, 
		output_MAC_1_30, output_MAC_1_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_2_0, output_MAC_2_1, output_MAC_2_2, output_MAC_2_3, output_MAC_2_4, output_MAC_2_5, output_MAC_2_6, output_MAC_2_7, output_MAC_2_8, output_MAC_2_9, 
		output_MAC_2_10, output_MAC_2_11, output_MAC_2_12, output_MAC_2_13, output_MAC_2_14, output_MAC_2_15, output_MAC_2_16, output_MAC_2_17, output_MAC_2_18, output_MAC_2_19, 
		output_MAC_2_20, output_MAC_2_21, output_MAC_2_22, output_MAC_2_23, output_MAC_2_24, output_MAC_2_25, output_MAC_2_26, output_MAC_2_27, output_MAC_2_28, output_MAC_2_29, 
		output_MAC_2_30, output_MAC_2_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_3_0, output_MAC_3_1, output_MAC_3_2, output_MAC_3_3, output_MAC_3_4, output_MAC_3_5, output_MAC_3_6, output_MAC_3_7, output_MAC_3_8, output_MAC_3_9, 
		output_MAC_3_10, output_MAC_3_11, output_MAC_3_12, output_MAC_3_13, output_MAC_3_14, output_MAC_3_15, output_MAC_3_16, output_MAC_3_17, output_MAC_3_18, output_MAC_3_19, 
		output_MAC_3_20, output_MAC_3_21, output_MAC_3_22, output_MAC_3_23, output_MAC_3_24, output_MAC_3_25, output_MAC_3_26, output_MAC_3_27, output_MAC_3_28, output_MAC_3_29, 
		output_MAC_3_30, output_MAC_3_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_4_0, output_MAC_4_1, output_MAC_4_2, output_MAC_4_3, output_MAC_4_4, output_MAC_4_5, output_MAC_4_6, output_MAC_4_7, output_MAC_4_8, output_MAC_4_9, 
		output_MAC_4_10, output_MAC_4_11, output_MAC_4_12, output_MAC_4_13, output_MAC_4_14, output_MAC_4_15, output_MAC_4_16, output_MAC_4_17, output_MAC_4_18, output_MAC_4_19, 
		output_MAC_4_20, output_MAC_4_21, output_MAC_4_22, output_MAC_4_23, output_MAC_4_24, output_MAC_4_25, output_MAC_4_26, output_MAC_4_27, output_MAC_4_28, output_MAC_4_29, 
		output_MAC_4_30, output_MAC_4_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_5_0, output_MAC_5_1, output_MAC_5_2, output_MAC_5_3, output_MAC_5_4, output_MAC_5_5, output_MAC_5_6, output_MAC_5_7, output_MAC_5_8, output_MAC_5_9, 
		output_MAC_5_10, output_MAC_5_11, output_MAC_5_12, output_MAC_5_13, output_MAC_5_14, output_MAC_5_15, output_MAC_5_16, output_MAC_5_17, output_MAC_5_18, output_MAC_5_19, 
		output_MAC_5_20, output_MAC_5_21, output_MAC_5_22, output_MAC_5_23, output_MAC_5_24, output_MAC_5_25, output_MAC_5_26, output_MAC_5_27, output_MAC_5_28, output_MAC_5_29, 
		output_MAC_5_30, output_MAC_5_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_6_0, output_MAC_6_1, output_MAC_6_2, output_MAC_6_3, output_MAC_6_4, output_MAC_6_5, output_MAC_6_6, output_MAC_6_7, output_MAC_6_8, output_MAC_6_9, 
		output_MAC_6_10, output_MAC_6_11, output_MAC_6_12, output_MAC_6_13, output_MAC_6_14, output_MAC_6_15, output_MAC_6_16, output_MAC_6_17, output_MAC_6_18, output_MAC_6_19, 
		output_MAC_6_20, output_MAC_6_21, output_MAC_6_22, output_MAC_6_23, output_MAC_6_24, output_MAC_6_25, output_MAC_6_26, output_MAC_6_27, output_MAC_6_28, output_MAC_6_29, 
		output_MAC_6_30, output_MAC_6_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_7_0, output_MAC_7_1, output_MAC_7_2, output_MAC_7_3, output_MAC_7_4, output_MAC_7_5, output_MAC_7_6, output_MAC_7_7, output_MAC_7_8, output_MAC_7_9, 
		output_MAC_7_10, output_MAC_7_11, output_MAC_7_12, output_MAC_7_13, output_MAC_7_14, output_MAC_7_15, output_MAC_7_16, output_MAC_7_17, output_MAC_7_18, output_MAC_7_19, 
		output_MAC_7_20, output_MAC_7_21, output_MAC_7_22, output_MAC_7_23, output_MAC_7_24, output_MAC_7_25, output_MAC_7_26, output_MAC_7_27, output_MAC_7_28, output_MAC_7_29, 
		output_MAC_7_30, output_MAC_7_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_8_0, output_MAC_8_1, output_MAC_8_2, output_MAC_8_3, output_MAC_8_4, output_MAC_8_5, output_MAC_8_6, output_MAC_8_7, output_MAC_8_8, output_MAC_8_9, 
		output_MAC_8_10, output_MAC_8_11, output_MAC_8_12, output_MAC_8_13, output_MAC_8_14, output_MAC_8_15, output_MAC_8_16, output_MAC_8_17, output_MAC_8_18, output_MAC_8_19, 
		output_MAC_8_20, output_MAC_8_21, output_MAC_8_22, output_MAC_8_23, output_MAC_8_24, output_MAC_8_25, output_MAC_8_26, output_MAC_8_27, output_MAC_8_28, output_MAC_8_29, 
		output_MAC_8_30, output_MAC_8_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_9_0, output_MAC_9_1, output_MAC_9_2, output_MAC_9_3, output_MAC_9_4, output_MAC_9_5, output_MAC_9_6, output_MAC_9_7, output_MAC_9_8, output_MAC_9_9, 
		output_MAC_9_10, output_MAC_9_11, output_MAC_9_12, output_MAC_9_13, output_MAC_9_14, output_MAC_9_15, output_MAC_9_16, output_MAC_9_17, output_MAC_9_18, output_MAC_9_19, 
		output_MAC_9_20, output_MAC_9_21, output_MAC_9_22, output_MAC_9_23, output_MAC_9_24, output_MAC_9_25, output_MAC_9_26, output_MAC_9_27, output_MAC_9_28, output_MAC_9_29, 
		output_MAC_9_30, output_MAC_9_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_10_0, output_MAC_10_1, output_MAC_10_2, output_MAC_10_3, output_MAC_10_4, output_MAC_10_5, output_MAC_10_6, output_MAC_10_7, output_MAC_10_8, output_MAC_10_9, 
		output_MAC_10_10, output_MAC_10_11, output_MAC_10_12, output_MAC_10_13, output_MAC_10_14, output_MAC_10_15, output_MAC_10_16, output_MAC_10_17, output_MAC_10_18, output_MAC_10_19, 
		output_MAC_10_20, output_MAC_10_21, output_MAC_10_22, output_MAC_10_23, output_MAC_10_24, output_MAC_10_25, output_MAC_10_26, output_MAC_10_27, output_MAC_10_28, output_MAC_10_29, 
		output_MAC_10_30, output_MAC_10_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_11_0, output_MAC_11_1, output_MAC_11_2, output_MAC_11_3, output_MAC_11_4, output_MAC_11_5, output_MAC_11_6, output_MAC_11_7, output_MAC_11_8, output_MAC_11_9, 
		output_MAC_11_10, output_MAC_11_11, output_MAC_11_12, output_MAC_11_13, output_MAC_11_14, output_MAC_11_15, output_MAC_11_16, output_MAC_11_17, output_MAC_11_18, output_MAC_11_19, 
		output_MAC_11_20, output_MAC_11_21, output_MAC_11_22, output_MAC_11_23, output_MAC_11_24, output_MAC_11_25, output_MAC_11_26, output_MAC_11_27, output_MAC_11_28, output_MAC_11_29, 
		output_MAC_11_30, output_MAC_11_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_12_0, output_MAC_12_1, output_MAC_12_2, output_MAC_12_3, output_MAC_12_4, output_MAC_12_5, output_MAC_12_6, output_MAC_12_7, output_MAC_12_8, output_MAC_12_9, 
		output_MAC_12_10, output_MAC_12_11, output_MAC_12_12, output_MAC_12_13, output_MAC_12_14, output_MAC_12_15, output_MAC_12_16, output_MAC_12_17, output_MAC_12_18, output_MAC_12_19, 
		output_MAC_12_20, output_MAC_12_21, output_MAC_12_22, output_MAC_12_23, output_MAC_12_24, output_MAC_12_25, output_MAC_12_26, output_MAC_12_27, output_MAC_12_28, output_MAC_12_29, 
		output_MAC_12_30, output_MAC_12_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_13_0, output_MAC_13_1, output_MAC_13_2, output_MAC_13_3, output_MAC_13_4, output_MAC_13_5, output_MAC_13_6, output_MAC_13_7, output_MAC_13_8, output_MAC_13_9, 
		output_MAC_13_10, output_MAC_13_11, output_MAC_13_12, output_MAC_13_13, output_MAC_13_14, output_MAC_13_15, output_MAC_13_16, output_MAC_13_17, output_MAC_13_18, output_MAC_13_19, 
		output_MAC_13_20, output_MAC_13_21, output_MAC_13_22, output_MAC_13_23, output_MAC_13_24, output_MAC_13_25, output_MAC_13_26, output_MAC_13_27, output_MAC_13_28, output_MAC_13_29, 
		output_MAC_13_30, output_MAC_13_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_14_0, output_MAC_14_1, output_MAC_14_2, output_MAC_14_3, output_MAC_14_4, output_MAC_14_5, output_MAC_14_6, output_MAC_14_7, output_MAC_14_8, output_MAC_14_9, 
		output_MAC_14_10, output_MAC_14_11, output_MAC_14_12, output_MAC_14_13, output_MAC_14_14, output_MAC_14_15, output_MAC_14_16, output_MAC_14_17, output_MAC_14_18, output_MAC_14_19, 
		output_MAC_14_20, output_MAC_14_21, output_MAC_14_22, output_MAC_14_23, output_MAC_14_24, output_MAC_14_25, output_MAC_14_26, output_MAC_14_27, output_MAC_14_28, output_MAC_14_29, 
		output_MAC_14_30, output_MAC_14_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_15_0, output_MAC_15_1, output_MAC_15_2, output_MAC_15_3, output_MAC_15_4, output_MAC_15_5, output_MAC_15_6, output_MAC_15_7, output_MAC_15_8, output_MAC_15_9, 
		output_MAC_15_10, output_MAC_15_11, output_MAC_15_12, output_MAC_15_13, output_MAC_15_14, output_MAC_15_15, output_MAC_15_16, output_MAC_15_17, output_MAC_15_18, output_MAC_15_19, 
		output_MAC_15_20, output_MAC_15_21, output_MAC_15_22, output_MAC_15_23, output_MAC_15_24, output_MAC_15_25, output_MAC_15_26, output_MAC_15_27, output_MAC_15_28, output_MAC_15_29, 
		output_MAC_15_30, output_MAC_15_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_16_0, output_MAC_16_1, output_MAC_16_2, output_MAC_16_3, output_MAC_16_4, output_MAC_16_5, output_MAC_16_6, output_MAC_16_7, output_MAC_16_8, output_MAC_16_9, 
		output_MAC_16_10, output_MAC_16_11, output_MAC_16_12, output_MAC_16_13, output_MAC_16_14, output_MAC_16_15, output_MAC_16_16, output_MAC_16_17, output_MAC_16_18, output_MAC_16_19, 
		output_MAC_16_20, output_MAC_16_21, output_MAC_16_22, output_MAC_16_23, output_MAC_16_24, output_MAC_16_25, output_MAC_16_26, output_MAC_16_27, output_MAC_16_28, output_MAC_16_29, 
		output_MAC_16_30, output_MAC_16_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_17_0, output_MAC_17_1, output_MAC_17_2, output_MAC_17_3, output_MAC_17_4, output_MAC_17_5, output_MAC_17_6, output_MAC_17_7, output_MAC_17_8, output_MAC_17_9, 
		output_MAC_17_10, output_MAC_17_11, output_MAC_17_12, output_MAC_17_13, output_MAC_17_14, output_MAC_17_15, output_MAC_17_16, output_MAC_17_17, output_MAC_17_18, output_MAC_17_19, 
		output_MAC_17_20, output_MAC_17_21, output_MAC_17_22, output_MAC_17_23, output_MAC_17_24, output_MAC_17_25, output_MAC_17_26, output_MAC_17_27, output_MAC_17_28, output_MAC_17_29, 
		output_MAC_17_30, output_MAC_17_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_18_0, output_MAC_18_1, output_MAC_18_2, output_MAC_18_3, output_MAC_18_4, output_MAC_18_5, output_MAC_18_6, output_MAC_18_7, output_MAC_18_8, output_MAC_18_9, 
		output_MAC_18_10, output_MAC_18_11, output_MAC_18_12, output_MAC_18_13, output_MAC_18_14, output_MAC_18_15, output_MAC_18_16, output_MAC_18_17, output_MAC_18_18, output_MAC_18_19, 
		output_MAC_18_20, output_MAC_18_21, output_MAC_18_22, output_MAC_18_23, output_MAC_18_24, output_MAC_18_25, output_MAC_18_26, output_MAC_18_27, output_MAC_18_28, output_MAC_18_29, 
		output_MAC_18_30, output_MAC_18_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_19_0, output_MAC_19_1, output_MAC_19_2, output_MAC_19_3, output_MAC_19_4, output_MAC_19_5, output_MAC_19_6, output_MAC_19_7, output_MAC_19_8, output_MAC_19_9, 
		output_MAC_19_10, output_MAC_19_11, output_MAC_19_12, output_MAC_19_13, output_MAC_19_14, output_MAC_19_15, output_MAC_19_16, output_MAC_19_17, output_MAC_19_18, output_MAC_19_19, 
		output_MAC_19_20, output_MAC_19_21, output_MAC_19_22, output_MAC_19_23, output_MAC_19_24, output_MAC_19_25, output_MAC_19_26, output_MAC_19_27, output_MAC_19_28, output_MAC_19_29, 
		output_MAC_19_30, output_MAC_19_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_20_0, output_MAC_20_1, output_MAC_20_2, output_MAC_20_3, output_MAC_20_4, output_MAC_20_5, output_MAC_20_6, output_MAC_20_7, output_MAC_20_8, output_MAC_20_9, 
		output_MAC_20_10, output_MAC_20_11, output_MAC_20_12, output_MAC_20_13, output_MAC_20_14, output_MAC_20_15, output_MAC_20_16, output_MAC_20_17, output_MAC_20_18, output_MAC_20_19, 
		output_MAC_20_20, output_MAC_20_21, output_MAC_20_22, output_MAC_20_23, output_MAC_20_24, output_MAC_20_25, output_MAC_20_26, output_MAC_20_27, output_MAC_20_28, output_MAC_20_29, 
		output_MAC_20_30, output_MAC_20_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_21_0, output_MAC_21_1, output_MAC_21_2, output_MAC_21_3, output_MAC_21_4, output_MAC_21_5, output_MAC_21_6, output_MAC_21_7, output_MAC_21_8, output_MAC_21_9, 
		output_MAC_21_10, output_MAC_21_11, output_MAC_21_12, output_MAC_21_13, output_MAC_21_14, output_MAC_21_15, output_MAC_21_16, output_MAC_21_17, output_MAC_21_18, output_MAC_21_19, 
		output_MAC_21_20, output_MAC_21_21, output_MAC_21_22, output_MAC_21_23, output_MAC_21_24, output_MAC_21_25, output_MAC_21_26, output_MAC_21_27, output_MAC_21_28, output_MAC_21_29, 
		output_MAC_21_30, output_MAC_21_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_22_0, output_MAC_22_1, output_MAC_22_2, output_MAC_22_3, output_MAC_22_4, output_MAC_22_5, output_MAC_22_6, output_MAC_22_7, output_MAC_22_8, output_MAC_22_9, 
		output_MAC_22_10, output_MAC_22_11, output_MAC_22_12, output_MAC_22_13, output_MAC_22_14, output_MAC_22_15, output_MAC_22_16, output_MAC_22_17, output_MAC_22_18, output_MAC_22_19, 
		output_MAC_22_20, output_MAC_22_21, output_MAC_22_22, output_MAC_22_23, output_MAC_22_24, output_MAC_22_25, output_MAC_22_26, output_MAC_22_27, output_MAC_22_28, output_MAC_22_29, 
		output_MAC_22_30, output_MAC_22_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_23_0, output_MAC_23_1, output_MAC_23_2, output_MAC_23_3, output_MAC_23_4, output_MAC_23_5, output_MAC_23_6, output_MAC_23_7, output_MAC_23_8, output_MAC_23_9, 
		output_MAC_23_10, output_MAC_23_11, output_MAC_23_12, output_MAC_23_13, output_MAC_23_14, output_MAC_23_15, output_MAC_23_16, output_MAC_23_17, output_MAC_23_18, output_MAC_23_19, 
		output_MAC_23_20, output_MAC_23_21, output_MAC_23_22, output_MAC_23_23, output_MAC_23_24, output_MAC_23_25, output_MAC_23_26, output_MAC_23_27, output_MAC_23_28, output_MAC_23_29, 
		output_MAC_23_30, output_MAC_23_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_24_0, output_MAC_24_1, output_MAC_24_2, output_MAC_24_3, output_MAC_24_4, output_MAC_24_5, output_MAC_24_6, output_MAC_24_7, output_MAC_24_8, output_MAC_24_9, 
		output_MAC_24_10, output_MAC_24_11, output_MAC_24_12, output_MAC_24_13, output_MAC_24_14, output_MAC_24_15, output_MAC_24_16, output_MAC_24_17, output_MAC_24_18, output_MAC_24_19, 
		output_MAC_24_20, output_MAC_24_21, output_MAC_24_22, output_MAC_24_23, output_MAC_24_24, output_MAC_24_25, output_MAC_24_26, output_MAC_24_27, output_MAC_24_28, output_MAC_24_29, 
		output_MAC_24_30, output_MAC_24_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_25_0, output_MAC_25_1, output_MAC_25_2, output_MAC_25_3, output_MAC_25_4, output_MAC_25_5, output_MAC_25_6, output_MAC_25_7, output_MAC_25_8, output_MAC_25_9, 
		output_MAC_25_10, output_MAC_25_11, output_MAC_25_12, output_MAC_25_13, output_MAC_25_14, output_MAC_25_15, output_MAC_25_16, output_MAC_25_17, output_MAC_25_18, output_MAC_25_19, 
		output_MAC_25_20, output_MAC_25_21, output_MAC_25_22, output_MAC_25_23, output_MAC_25_24, output_MAC_25_25, output_MAC_25_26, output_MAC_25_27, output_MAC_25_28, output_MAC_25_29, 
		output_MAC_25_30, output_MAC_25_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_26_0, output_MAC_26_1, output_MAC_26_2, output_MAC_26_3, output_MAC_26_4, output_MAC_26_5, output_MAC_26_6, output_MAC_26_7, output_MAC_26_8, output_MAC_26_9, 
		output_MAC_26_10, output_MAC_26_11, output_MAC_26_12, output_MAC_26_13, output_MAC_26_14, output_MAC_26_15, output_MAC_26_16, output_MAC_26_17, output_MAC_26_18, output_MAC_26_19, 
		output_MAC_26_20, output_MAC_26_21, output_MAC_26_22, output_MAC_26_23, output_MAC_26_24, output_MAC_26_25, output_MAC_26_26, output_MAC_26_27, output_MAC_26_28, output_MAC_26_29, 
		output_MAC_26_30, output_MAC_26_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_27_0, output_MAC_27_1, output_MAC_27_2, output_MAC_27_3, output_MAC_27_4, output_MAC_27_5, output_MAC_27_6, output_MAC_27_7, output_MAC_27_8, output_MAC_27_9, 
		output_MAC_27_10, output_MAC_27_11, output_MAC_27_12, output_MAC_27_13, output_MAC_27_14, output_MAC_27_15, output_MAC_27_16, output_MAC_27_17, output_MAC_27_18, output_MAC_27_19, 
		output_MAC_27_20, output_MAC_27_21, output_MAC_27_22, output_MAC_27_23, output_MAC_27_24, output_MAC_27_25, output_MAC_27_26, output_MAC_27_27, output_MAC_27_28, output_MAC_27_29, 
		output_MAC_27_30, output_MAC_27_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_28_0, output_MAC_28_1, output_MAC_28_2, output_MAC_28_3, output_MAC_28_4, output_MAC_28_5, output_MAC_28_6, output_MAC_28_7, output_MAC_28_8, output_MAC_28_9, 
		output_MAC_28_10, output_MAC_28_11, output_MAC_28_12, output_MAC_28_13, output_MAC_28_14, output_MAC_28_15, output_MAC_28_16, output_MAC_28_17, output_MAC_28_18, output_MAC_28_19, 
		output_MAC_28_20, output_MAC_28_21, output_MAC_28_22, output_MAC_28_23, output_MAC_28_24, output_MAC_28_25, output_MAC_28_26, output_MAC_28_27, output_MAC_28_28, output_MAC_28_29, 
		output_MAC_28_30, output_MAC_28_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_29_0, output_MAC_29_1, output_MAC_29_2, output_MAC_29_3, output_MAC_29_4, output_MAC_29_5, output_MAC_29_6, output_MAC_29_7, output_MAC_29_8, output_MAC_29_9, 
		output_MAC_29_10, output_MAC_29_11, output_MAC_29_12, output_MAC_29_13, output_MAC_29_14, output_MAC_29_15, output_MAC_29_16, output_MAC_29_17, output_MAC_29_18, output_MAC_29_19, 
		output_MAC_29_20, output_MAC_29_21, output_MAC_29_22, output_MAC_29_23, output_MAC_29_24, output_MAC_29_25, output_MAC_29_26, output_MAC_29_27, output_MAC_29_28, output_MAC_29_29, 
		output_MAC_29_30, output_MAC_29_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_30_0, output_MAC_30_1, output_MAC_30_2, output_MAC_30_3, output_MAC_30_4, output_MAC_30_5, output_MAC_30_6, output_MAC_30_7, output_MAC_30_8, output_MAC_30_9, 
		output_MAC_30_10, output_MAC_30_11, output_MAC_30_12, output_MAC_30_13, output_MAC_30_14, output_MAC_30_15, output_MAC_30_16, output_MAC_30_17, output_MAC_30_18, output_MAC_30_19, 
		output_MAC_30_20, output_MAC_30_21, output_MAC_30_22, output_MAC_30_23, output_MAC_30_24, output_MAC_30_25, output_MAC_30_26, output_MAC_30_27, output_MAC_30_28, output_MAC_30_29, 
		output_MAC_30_30, output_MAC_30_31: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_31_0, output_MAC_31_1, output_MAC_31_2, output_MAC_31_3, output_MAC_31_4, output_MAC_31_5, output_MAC_31_6, output_MAC_31_7, output_MAC_31_8, output_MAC_31_9, 
		output_MAC_31_10, output_MAC_31_11, output_MAC_31_12, output_MAC_31_13, output_MAC_31_14, output_MAC_31_15, output_MAC_31_16, output_MAC_31_17, output_MAC_31_18, output_MAC_31_19, 
		output_MAC_31_20, output_MAC_31_21, output_MAC_31_22, output_MAC_31_23, output_MAC_31_24, output_MAC_31_25, output_MAC_31_26, output_MAC_31_27, output_MAC_31_28, output_MAC_31_29, 
		output_MAC_31_30, output_MAC_31_31: STD_LOGIC_VECTOR(31 downto 0);

BEGIN

	input_row_0_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_0, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_0);
	input_row_1_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_1, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_1);
	input_row_2_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_2, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_2);
	input_row_3_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_3, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_3);
	input_row_4_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_4, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_4);
	input_row_5_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_5, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_5);
	input_row_6_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_6, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_6);
	input_row_7_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_7, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_7);
	input_row_8_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_8, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_8);
	input_row_9_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_9, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_9);
	input_row_10_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_10, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_10);
	input_row_11_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_11, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_11);
	input_row_12_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_12, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_12);
	input_row_13_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_13, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_13);
	input_row_14_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_14, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_14);
	input_row_15_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_15, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_15);
	input_row_16_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_16, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_16);
	input_row_17_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_17, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_17);
	input_row_18_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_18, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_18);
	input_row_19_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_19, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_19);
	input_row_20_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_20, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_20);
	input_row_21_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_21, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_21);
	input_row_22_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_22, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_22);
	input_row_23_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_23, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_23);
	input_row_24_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_24, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_24);
	input_row_25_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_25, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_25);
	input_row_26_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_26, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_26);
	input_row_27_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_27, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_27);
	input_row_28_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_28, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_28);
	input_row_29_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_29, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_29);
	input_row_30_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_30, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_30);
	input_row_31_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_row_31, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_row_31);
	input_col_0_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_0, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_0);

	input_col_1_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_1, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_1);

	input_col_2_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_2, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_2);

	input_col_3_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_3, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_3);

	input_col_4_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_4, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_4);

	input_col_5_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_5, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_5);

	input_col_6_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_6, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_6);

	input_col_7_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_7, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_7);

	input_col_8_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_8, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_8);

	input_col_9_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_9, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_9);

	input_col_10_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_10, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_10);

	input_col_11_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_11, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_11);

	input_col_12_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_12, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_12);

	input_col_13_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_13, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_13);

	input_col_14_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_14, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_14);

	input_col_15_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_15, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_15);

	input_col_16_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_16, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_16);

	input_col_17_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_17, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_17);

	input_col_18_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_18, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_18);

	input_col_19_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_19, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_19);

	input_col_20_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_20, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_20);

	input_col_21_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_21, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_21);

	input_col_22_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_22, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_22);

	input_col_23_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_23, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_23);

	input_col_24_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_24, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_24);

	input_col_25_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_25, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_25);

	input_col_26_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_26, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_26);

	input_col_27_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_27, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_27);

	input_col_28_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_28, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_28);

	input_col_29_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_29, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_29);

	input_col_30_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_30, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_30);

	input_col_31_reg: regnbit GENERIC MAP(N=>8)
		PORT MAP(D=>input_col_31, CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, Q=>reg_input_col_31);

	enable_ff_in: ff PORT MAP(D=>ENABLE, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>reg_ENABLE_in);
	sel_mux_reg: regnbit GENERIC MAP(N=>5) PORT MAP(D=>SEL_MUX, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>reg_SEL_MUX);

	MAC_0_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_0, data_out=>output_MAC_0_0);

	MAC_0_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_1, data_out=>output_MAC_0_1);

	MAC_0_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_2, data_out=>output_MAC_0_2);

	MAC_0_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_3, data_out=>output_MAC_0_3);

	MAC_0_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_4, data_out=>output_MAC_0_4);

	MAC_0_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_5, data_out=>output_MAC_0_5);

	MAC_0_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_6, data_out=>output_MAC_0_6);

	MAC_0_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_7, data_out=>output_MAC_0_7);

	MAC_0_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_8, data_out=>output_MAC_0_8);

	MAC_0_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_9, data_out=>output_MAC_0_9);

	MAC_0_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_10, data_out=>output_MAC_0_10);

	MAC_0_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_11, data_out=>output_MAC_0_11);

	MAC_0_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_12, data_out=>output_MAC_0_12);

	MAC_0_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_13, data_out=>output_MAC_0_13);

	MAC_0_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_14, data_out=>output_MAC_0_14);

	MAC_0_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_15, data_out=>output_MAC_0_15);

	MAC_0_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_16, data_out=>output_MAC_0_16);

	MAC_0_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_17, data_out=>output_MAC_0_17);

	MAC_0_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_18, data_out=>output_MAC_0_18);

	MAC_0_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_19, data_out=>output_MAC_0_19);

	MAC_0_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_20, data_out=>output_MAC_0_20);

	MAC_0_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_21, data_out=>output_MAC_0_21);

	MAC_0_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_22, data_out=>output_MAC_0_22);

	MAC_0_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_23, data_out=>output_MAC_0_23);

	MAC_0_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_24, data_out=>output_MAC_0_24);

	MAC_0_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_25, data_out=>output_MAC_0_25);

	MAC_0_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_26, data_out=>output_MAC_0_26);

	MAC_0_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_27, data_out=>output_MAC_0_27);

	MAC_0_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_28, data_out=>output_MAC_0_28);

	MAC_0_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_29, data_out=>output_MAC_0_29);

	MAC_0_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_30, data_out=>output_MAC_0_30);

	MAC_0_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_0, data_in_B=>reg_input_col_31, data_out=>output_MAC_0_31);

	MAC_1_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_0, data_out=>output_MAC_1_0);

	MAC_1_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_1, data_out=>output_MAC_1_1);

	MAC_1_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_2, data_out=>output_MAC_1_2);

	MAC_1_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_3, data_out=>output_MAC_1_3);

	MAC_1_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_4, data_out=>output_MAC_1_4);

	MAC_1_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_5, data_out=>output_MAC_1_5);

	MAC_1_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_6, data_out=>output_MAC_1_6);

	MAC_1_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_7, data_out=>output_MAC_1_7);

	MAC_1_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_8, data_out=>output_MAC_1_8);

	MAC_1_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_9, data_out=>output_MAC_1_9);

	MAC_1_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_10, data_out=>output_MAC_1_10);

	MAC_1_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_11, data_out=>output_MAC_1_11);

	MAC_1_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_12, data_out=>output_MAC_1_12);

	MAC_1_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_13, data_out=>output_MAC_1_13);

	MAC_1_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_14, data_out=>output_MAC_1_14);

	MAC_1_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_15, data_out=>output_MAC_1_15);

	MAC_1_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_16, data_out=>output_MAC_1_16);

	MAC_1_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_17, data_out=>output_MAC_1_17);

	MAC_1_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_18, data_out=>output_MAC_1_18);

	MAC_1_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_19, data_out=>output_MAC_1_19);

	MAC_1_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_20, data_out=>output_MAC_1_20);

	MAC_1_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_21, data_out=>output_MAC_1_21);

	MAC_1_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_22, data_out=>output_MAC_1_22);

	MAC_1_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_23, data_out=>output_MAC_1_23);

	MAC_1_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_24, data_out=>output_MAC_1_24);

	MAC_1_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_25, data_out=>output_MAC_1_25);

	MAC_1_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_26, data_out=>output_MAC_1_26);

	MAC_1_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_27, data_out=>output_MAC_1_27);

	MAC_1_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_28, data_out=>output_MAC_1_28);

	MAC_1_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_29, data_out=>output_MAC_1_29);

	MAC_1_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_30, data_out=>output_MAC_1_30);

	MAC_1_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_1, data_in_B=>reg_input_col_31, data_out=>output_MAC_1_31);

	MAC_2_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_0, data_out=>output_MAC_2_0);

	MAC_2_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_1, data_out=>output_MAC_2_1);

	MAC_2_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_2, data_out=>output_MAC_2_2);

	MAC_2_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_3, data_out=>output_MAC_2_3);

	MAC_2_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_4, data_out=>output_MAC_2_4);

	MAC_2_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_5, data_out=>output_MAC_2_5);

	MAC_2_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_6, data_out=>output_MAC_2_6);

	MAC_2_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_7, data_out=>output_MAC_2_7);

	MAC_2_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_8, data_out=>output_MAC_2_8);

	MAC_2_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_9, data_out=>output_MAC_2_9);

	MAC_2_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_10, data_out=>output_MAC_2_10);

	MAC_2_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_11, data_out=>output_MAC_2_11);

	MAC_2_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_12, data_out=>output_MAC_2_12);

	MAC_2_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_13, data_out=>output_MAC_2_13);

	MAC_2_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_14, data_out=>output_MAC_2_14);

	MAC_2_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_15, data_out=>output_MAC_2_15);

	MAC_2_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_16, data_out=>output_MAC_2_16);

	MAC_2_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_17, data_out=>output_MAC_2_17);

	MAC_2_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_18, data_out=>output_MAC_2_18);

	MAC_2_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_19, data_out=>output_MAC_2_19);

	MAC_2_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_20, data_out=>output_MAC_2_20);

	MAC_2_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_21, data_out=>output_MAC_2_21);

	MAC_2_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_22, data_out=>output_MAC_2_22);

	MAC_2_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_23, data_out=>output_MAC_2_23);

	MAC_2_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_24, data_out=>output_MAC_2_24);

	MAC_2_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_25, data_out=>output_MAC_2_25);

	MAC_2_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_26, data_out=>output_MAC_2_26);

	MAC_2_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_27, data_out=>output_MAC_2_27);

	MAC_2_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_28, data_out=>output_MAC_2_28);

	MAC_2_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_29, data_out=>output_MAC_2_29);

	MAC_2_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_30, data_out=>output_MAC_2_30);

	MAC_2_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_2, data_in_B=>reg_input_col_31, data_out=>output_MAC_2_31);

	MAC_3_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_0, data_out=>output_MAC_3_0);

	MAC_3_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_1, data_out=>output_MAC_3_1);

	MAC_3_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_2, data_out=>output_MAC_3_2);

	MAC_3_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_3, data_out=>output_MAC_3_3);

	MAC_3_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_4, data_out=>output_MAC_3_4);

	MAC_3_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_5, data_out=>output_MAC_3_5);

	MAC_3_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_6, data_out=>output_MAC_3_6);

	MAC_3_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_7, data_out=>output_MAC_3_7);

	MAC_3_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_8, data_out=>output_MAC_3_8);

	MAC_3_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_9, data_out=>output_MAC_3_9);

	MAC_3_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_10, data_out=>output_MAC_3_10);

	MAC_3_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_11, data_out=>output_MAC_3_11);

	MAC_3_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_12, data_out=>output_MAC_3_12);

	MAC_3_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_13, data_out=>output_MAC_3_13);

	MAC_3_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_14, data_out=>output_MAC_3_14);

	MAC_3_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_15, data_out=>output_MAC_3_15);

	MAC_3_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_16, data_out=>output_MAC_3_16);

	MAC_3_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_17, data_out=>output_MAC_3_17);

	MAC_3_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_18, data_out=>output_MAC_3_18);

	MAC_3_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_19, data_out=>output_MAC_3_19);

	MAC_3_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_20, data_out=>output_MAC_3_20);

	MAC_3_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_21, data_out=>output_MAC_3_21);

	MAC_3_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_22, data_out=>output_MAC_3_22);

	MAC_3_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_23, data_out=>output_MAC_3_23);

	MAC_3_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_24, data_out=>output_MAC_3_24);

	MAC_3_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_25, data_out=>output_MAC_3_25);

	MAC_3_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_26, data_out=>output_MAC_3_26);

	MAC_3_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_27, data_out=>output_MAC_3_27);

	MAC_3_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_28, data_out=>output_MAC_3_28);

	MAC_3_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_29, data_out=>output_MAC_3_29);

	MAC_3_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_30, data_out=>output_MAC_3_30);

	MAC_3_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_3, data_in_B=>reg_input_col_31, data_out=>output_MAC_3_31);

	MAC_4_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_0, data_out=>output_MAC_4_0);

	MAC_4_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_1, data_out=>output_MAC_4_1);

	MAC_4_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_2, data_out=>output_MAC_4_2);

	MAC_4_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_3, data_out=>output_MAC_4_3);

	MAC_4_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_4, data_out=>output_MAC_4_4);

	MAC_4_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_5, data_out=>output_MAC_4_5);

	MAC_4_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_6, data_out=>output_MAC_4_6);

	MAC_4_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_7, data_out=>output_MAC_4_7);

	MAC_4_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_8, data_out=>output_MAC_4_8);

	MAC_4_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_9, data_out=>output_MAC_4_9);

	MAC_4_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_10, data_out=>output_MAC_4_10);

	MAC_4_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_11, data_out=>output_MAC_4_11);

	MAC_4_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_12, data_out=>output_MAC_4_12);

	MAC_4_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_13, data_out=>output_MAC_4_13);

	MAC_4_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_14, data_out=>output_MAC_4_14);

	MAC_4_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_15, data_out=>output_MAC_4_15);

	MAC_4_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_16, data_out=>output_MAC_4_16);

	MAC_4_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_17, data_out=>output_MAC_4_17);

	MAC_4_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_18, data_out=>output_MAC_4_18);

	MAC_4_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_19, data_out=>output_MAC_4_19);

	MAC_4_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_20, data_out=>output_MAC_4_20);

	MAC_4_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_21, data_out=>output_MAC_4_21);

	MAC_4_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_22, data_out=>output_MAC_4_22);

	MAC_4_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_23, data_out=>output_MAC_4_23);

	MAC_4_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_24, data_out=>output_MAC_4_24);

	MAC_4_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_25, data_out=>output_MAC_4_25);

	MAC_4_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_26, data_out=>output_MAC_4_26);

	MAC_4_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_27, data_out=>output_MAC_4_27);

	MAC_4_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_28, data_out=>output_MAC_4_28);

	MAC_4_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_29, data_out=>output_MAC_4_29);

	MAC_4_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_30, data_out=>output_MAC_4_30);

	MAC_4_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_4, data_in_B=>reg_input_col_31, data_out=>output_MAC_4_31);

	MAC_5_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_0, data_out=>output_MAC_5_0);

	MAC_5_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_1, data_out=>output_MAC_5_1);

	MAC_5_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_2, data_out=>output_MAC_5_2);

	MAC_5_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_3, data_out=>output_MAC_5_3);

	MAC_5_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_4, data_out=>output_MAC_5_4);

	MAC_5_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_5, data_out=>output_MAC_5_5);

	MAC_5_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_6, data_out=>output_MAC_5_6);

	MAC_5_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_7, data_out=>output_MAC_5_7);

	MAC_5_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_8, data_out=>output_MAC_5_8);

	MAC_5_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_9, data_out=>output_MAC_5_9);

	MAC_5_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_10, data_out=>output_MAC_5_10);

	MAC_5_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_11, data_out=>output_MAC_5_11);

	MAC_5_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_12, data_out=>output_MAC_5_12);

	MAC_5_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_13, data_out=>output_MAC_5_13);

	MAC_5_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_14, data_out=>output_MAC_5_14);

	MAC_5_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_15, data_out=>output_MAC_5_15);

	MAC_5_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_16, data_out=>output_MAC_5_16);

	MAC_5_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_17, data_out=>output_MAC_5_17);

	MAC_5_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_18, data_out=>output_MAC_5_18);

	MAC_5_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_19, data_out=>output_MAC_5_19);

	MAC_5_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_20, data_out=>output_MAC_5_20);

	MAC_5_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_21, data_out=>output_MAC_5_21);

	MAC_5_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_22, data_out=>output_MAC_5_22);

	MAC_5_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_23, data_out=>output_MAC_5_23);

	MAC_5_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_24, data_out=>output_MAC_5_24);

	MAC_5_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_25, data_out=>output_MAC_5_25);

	MAC_5_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_26, data_out=>output_MAC_5_26);

	MAC_5_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_27, data_out=>output_MAC_5_27);

	MAC_5_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_28, data_out=>output_MAC_5_28);

	MAC_5_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_29, data_out=>output_MAC_5_29);

	MAC_5_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_30, data_out=>output_MAC_5_30);

	MAC_5_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_5, data_in_B=>reg_input_col_31, data_out=>output_MAC_5_31);

	MAC_6_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_0, data_out=>output_MAC_6_0);

	MAC_6_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_1, data_out=>output_MAC_6_1);

	MAC_6_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_2, data_out=>output_MAC_6_2);

	MAC_6_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_3, data_out=>output_MAC_6_3);

	MAC_6_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_4, data_out=>output_MAC_6_4);

	MAC_6_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_5, data_out=>output_MAC_6_5);

	MAC_6_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_6, data_out=>output_MAC_6_6);

	MAC_6_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_7, data_out=>output_MAC_6_7);

	MAC_6_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_8, data_out=>output_MAC_6_8);

	MAC_6_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_9, data_out=>output_MAC_6_9);

	MAC_6_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_10, data_out=>output_MAC_6_10);

	MAC_6_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_11, data_out=>output_MAC_6_11);

	MAC_6_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_12, data_out=>output_MAC_6_12);

	MAC_6_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_13, data_out=>output_MAC_6_13);

	MAC_6_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_14, data_out=>output_MAC_6_14);

	MAC_6_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_15, data_out=>output_MAC_6_15);

	MAC_6_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_16, data_out=>output_MAC_6_16);

	MAC_6_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_17, data_out=>output_MAC_6_17);

	MAC_6_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_18, data_out=>output_MAC_6_18);

	MAC_6_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_19, data_out=>output_MAC_6_19);

	MAC_6_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_20, data_out=>output_MAC_6_20);

	MAC_6_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_21, data_out=>output_MAC_6_21);

	MAC_6_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_22, data_out=>output_MAC_6_22);

	MAC_6_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_23, data_out=>output_MAC_6_23);

	MAC_6_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_24, data_out=>output_MAC_6_24);

	MAC_6_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_25, data_out=>output_MAC_6_25);

	MAC_6_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_26, data_out=>output_MAC_6_26);

	MAC_6_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_27, data_out=>output_MAC_6_27);

	MAC_6_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_28, data_out=>output_MAC_6_28);

	MAC_6_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_29, data_out=>output_MAC_6_29);

	MAC_6_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_30, data_out=>output_MAC_6_30);

	MAC_6_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_6, data_in_B=>reg_input_col_31, data_out=>output_MAC_6_31);

	MAC_7_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_0, data_out=>output_MAC_7_0);

	MAC_7_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_1, data_out=>output_MAC_7_1);

	MAC_7_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_2, data_out=>output_MAC_7_2);

	MAC_7_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_3, data_out=>output_MAC_7_3);

	MAC_7_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_4, data_out=>output_MAC_7_4);

	MAC_7_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_5, data_out=>output_MAC_7_5);

	MAC_7_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_6, data_out=>output_MAC_7_6);

	MAC_7_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_7, data_out=>output_MAC_7_7);

	MAC_7_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_8, data_out=>output_MAC_7_8);

	MAC_7_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_9, data_out=>output_MAC_7_9);

	MAC_7_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_10, data_out=>output_MAC_7_10);

	MAC_7_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_11, data_out=>output_MAC_7_11);

	MAC_7_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_12, data_out=>output_MAC_7_12);

	MAC_7_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_13, data_out=>output_MAC_7_13);

	MAC_7_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_14, data_out=>output_MAC_7_14);

	MAC_7_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_15, data_out=>output_MAC_7_15);

	MAC_7_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_16, data_out=>output_MAC_7_16);

	MAC_7_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_17, data_out=>output_MAC_7_17);

	MAC_7_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_18, data_out=>output_MAC_7_18);

	MAC_7_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_19, data_out=>output_MAC_7_19);

	MAC_7_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_20, data_out=>output_MAC_7_20);

	MAC_7_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_21, data_out=>output_MAC_7_21);

	MAC_7_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_22, data_out=>output_MAC_7_22);

	MAC_7_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_23, data_out=>output_MAC_7_23);

	MAC_7_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_24, data_out=>output_MAC_7_24);

	MAC_7_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_25, data_out=>output_MAC_7_25);

	MAC_7_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_26, data_out=>output_MAC_7_26);

	MAC_7_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_27, data_out=>output_MAC_7_27);

	MAC_7_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_28, data_out=>output_MAC_7_28);

	MAC_7_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_29, data_out=>output_MAC_7_29);

	MAC_7_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_30, data_out=>output_MAC_7_30);

	MAC_7_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_7, data_in_B=>reg_input_col_31, data_out=>output_MAC_7_31);

	MAC_8_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_0, data_out=>output_MAC_8_0);

	MAC_8_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_1, data_out=>output_MAC_8_1);

	MAC_8_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_2, data_out=>output_MAC_8_2);

	MAC_8_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_3, data_out=>output_MAC_8_3);

	MAC_8_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_4, data_out=>output_MAC_8_4);

	MAC_8_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_5, data_out=>output_MAC_8_5);

	MAC_8_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_6, data_out=>output_MAC_8_6);

	MAC_8_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_7, data_out=>output_MAC_8_7);

	MAC_8_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_8, data_out=>output_MAC_8_8);

	MAC_8_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_9, data_out=>output_MAC_8_9);

	MAC_8_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_10, data_out=>output_MAC_8_10);

	MAC_8_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_11, data_out=>output_MAC_8_11);

	MAC_8_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_12, data_out=>output_MAC_8_12);

	MAC_8_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_13, data_out=>output_MAC_8_13);

	MAC_8_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_14, data_out=>output_MAC_8_14);

	MAC_8_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_15, data_out=>output_MAC_8_15);

	MAC_8_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_16, data_out=>output_MAC_8_16);

	MAC_8_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_17, data_out=>output_MAC_8_17);

	MAC_8_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_18, data_out=>output_MAC_8_18);

	MAC_8_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_19, data_out=>output_MAC_8_19);

	MAC_8_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_20, data_out=>output_MAC_8_20);

	MAC_8_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_21, data_out=>output_MAC_8_21);

	MAC_8_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_22, data_out=>output_MAC_8_22);

	MAC_8_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_23, data_out=>output_MAC_8_23);

	MAC_8_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_24, data_out=>output_MAC_8_24);

	MAC_8_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_25, data_out=>output_MAC_8_25);

	MAC_8_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_26, data_out=>output_MAC_8_26);

	MAC_8_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_27, data_out=>output_MAC_8_27);

	MAC_8_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_28, data_out=>output_MAC_8_28);

	MAC_8_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_29, data_out=>output_MAC_8_29);

	MAC_8_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_30, data_out=>output_MAC_8_30);

	MAC_8_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_8, data_in_B=>reg_input_col_31, data_out=>output_MAC_8_31);

	MAC_9_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_0, data_out=>output_MAC_9_0);

	MAC_9_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_1, data_out=>output_MAC_9_1);

	MAC_9_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_2, data_out=>output_MAC_9_2);

	MAC_9_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_3, data_out=>output_MAC_9_3);

	MAC_9_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_4, data_out=>output_MAC_9_4);

	MAC_9_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_5, data_out=>output_MAC_9_5);

	MAC_9_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_6, data_out=>output_MAC_9_6);

	MAC_9_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_7, data_out=>output_MAC_9_7);

	MAC_9_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_8, data_out=>output_MAC_9_8);

	MAC_9_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_9, data_out=>output_MAC_9_9);

	MAC_9_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_10, data_out=>output_MAC_9_10);

	MAC_9_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_11, data_out=>output_MAC_9_11);

	MAC_9_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_12, data_out=>output_MAC_9_12);

	MAC_9_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_13, data_out=>output_MAC_9_13);

	MAC_9_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_14, data_out=>output_MAC_9_14);

	MAC_9_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_15, data_out=>output_MAC_9_15);

	MAC_9_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_16, data_out=>output_MAC_9_16);

	MAC_9_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_17, data_out=>output_MAC_9_17);

	MAC_9_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_18, data_out=>output_MAC_9_18);

	MAC_9_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_19, data_out=>output_MAC_9_19);

	MAC_9_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_20, data_out=>output_MAC_9_20);

	MAC_9_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_21, data_out=>output_MAC_9_21);

	MAC_9_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_22, data_out=>output_MAC_9_22);

	MAC_9_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_23, data_out=>output_MAC_9_23);

	MAC_9_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_24, data_out=>output_MAC_9_24);

	MAC_9_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_25, data_out=>output_MAC_9_25);

	MAC_9_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_26, data_out=>output_MAC_9_26);

	MAC_9_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_27, data_out=>output_MAC_9_27);

	MAC_9_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_28, data_out=>output_MAC_9_28);

	MAC_9_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_29, data_out=>output_MAC_9_29);

	MAC_9_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_30, data_out=>output_MAC_9_30);

	MAC_9_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_9, data_in_B=>reg_input_col_31, data_out=>output_MAC_9_31);

	MAC_10_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_0, data_out=>output_MAC_10_0);

	MAC_10_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_1, data_out=>output_MAC_10_1);

	MAC_10_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_2, data_out=>output_MAC_10_2);

	MAC_10_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_3, data_out=>output_MAC_10_3);

	MAC_10_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_4, data_out=>output_MAC_10_4);

	MAC_10_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_5, data_out=>output_MAC_10_5);

	MAC_10_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_6, data_out=>output_MAC_10_6);

	MAC_10_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_7, data_out=>output_MAC_10_7);

	MAC_10_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_8, data_out=>output_MAC_10_8);

	MAC_10_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_9, data_out=>output_MAC_10_9);

	MAC_10_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_10, data_out=>output_MAC_10_10);

	MAC_10_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_11, data_out=>output_MAC_10_11);

	MAC_10_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_12, data_out=>output_MAC_10_12);

	MAC_10_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_13, data_out=>output_MAC_10_13);

	MAC_10_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_14, data_out=>output_MAC_10_14);

	MAC_10_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_15, data_out=>output_MAC_10_15);

	MAC_10_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_16, data_out=>output_MAC_10_16);

	MAC_10_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_17, data_out=>output_MAC_10_17);

	MAC_10_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_18, data_out=>output_MAC_10_18);

	MAC_10_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_19, data_out=>output_MAC_10_19);

	MAC_10_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_20, data_out=>output_MAC_10_20);

	MAC_10_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_21, data_out=>output_MAC_10_21);

	MAC_10_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_22, data_out=>output_MAC_10_22);

	MAC_10_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_23, data_out=>output_MAC_10_23);

	MAC_10_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_24, data_out=>output_MAC_10_24);

	MAC_10_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_25, data_out=>output_MAC_10_25);

	MAC_10_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_26, data_out=>output_MAC_10_26);

	MAC_10_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_27, data_out=>output_MAC_10_27);

	MAC_10_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_28, data_out=>output_MAC_10_28);

	MAC_10_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_29, data_out=>output_MAC_10_29);

	MAC_10_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_30, data_out=>output_MAC_10_30);

	MAC_10_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_10, data_in_B=>reg_input_col_31, data_out=>output_MAC_10_31);

	MAC_11_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_0, data_out=>output_MAC_11_0);

	MAC_11_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_1, data_out=>output_MAC_11_1);

	MAC_11_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_2, data_out=>output_MAC_11_2);

	MAC_11_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_3, data_out=>output_MAC_11_3);

	MAC_11_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_4, data_out=>output_MAC_11_4);

	MAC_11_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_5, data_out=>output_MAC_11_5);

	MAC_11_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_6, data_out=>output_MAC_11_6);

	MAC_11_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_7, data_out=>output_MAC_11_7);

	MAC_11_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_8, data_out=>output_MAC_11_8);

	MAC_11_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_9, data_out=>output_MAC_11_9);

	MAC_11_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_10, data_out=>output_MAC_11_10);

	MAC_11_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_11, data_out=>output_MAC_11_11);

	MAC_11_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_12, data_out=>output_MAC_11_12);

	MAC_11_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_13, data_out=>output_MAC_11_13);

	MAC_11_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_14, data_out=>output_MAC_11_14);

	MAC_11_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_15, data_out=>output_MAC_11_15);

	MAC_11_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_16, data_out=>output_MAC_11_16);

	MAC_11_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_17, data_out=>output_MAC_11_17);

	MAC_11_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_18, data_out=>output_MAC_11_18);

	MAC_11_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_19, data_out=>output_MAC_11_19);

	MAC_11_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_20, data_out=>output_MAC_11_20);

	MAC_11_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_21, data_out=>output_MAC_11_21);

	MAC_11_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_22, data_out=>output_MAC_11_22);

	MAC_11_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_23, data_out=>output_MAC_11_23);

	MAC_11_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_24, data_out=>output_MAC_11_24);

	MAC_11_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_25, data_out=>output_MAC_11_25);

	MAC_11_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_26, data_out=>output_MAC_11_26);

	MAC_11_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_27, data_out=>output_MAC_11_27);

	MAC_11_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_28, data_out=>output_MAC_11_28);

	MAC_11_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_29, data_out=>output_MAC_11_29);

	MAC_11_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_30, data_out=>output_MAC_11_30);

	MAC_11_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_11, data_in_B=>reg_input_col_31, data_out=>output_MAC_11_31);

	MAC_12_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_0, data_out=>output_MAC_12_0);

	MAC_12_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_1, data_out=>output_MAC_12_1);

	MAC_12_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_2, data_out=>output_MAC_12_2);

	MAC_12_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_3, data_out=>output_MAC_12_3);

	MAC_12_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_4, data_out=>output_MAC_12_4);

	MAC_12_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_5, data_out=>output_MAC_12_5);

	MAC_12_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_6, data_out=>output_MAC_12_6);

	MAC_12_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_7, data_out=>output_MAC_12_7);

	MAC_12_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_8, data_out=>output_MAC_12_8);

	MAC_12_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_9, data_out=>output_MAC_12_9);

	MAC_12_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_10, data_out=>output_MAC_12_10);

	MAC_12_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_11, data_out=>output_MAC_12_11);

	MAC_12_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_12, data_out=>output_MAC_12_12);

	MAC_12_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_13, data_out=>output_MAC_12_13);

	MAC_12_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_14, data_out=>output_MAC_12_14);

	MAC_12_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_15, data_out=>output_MAC_12_15);

	MAC_12_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_16, data_out=>output_MAC_12_16);

	MAC_12_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_17, data_out=>output_MAC_12_17);

	MAC_12_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_18, data_out=>output_MAC_12_18);

	MAC_12_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_19, data_out=>output_MAC_12_19);

	MAC_12_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_20, data_out=>output_MAC_12_20);

	MAC_12_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_21, data_out=>output_MAC_12_21);

	MAC_12_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_22, data_out=>output_MAC_12_22);

	MAC_12_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_23, data_out=>output_MAC_12_23);

	MAC_12_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_24, data_out=>output_MAC_12_24);

	MAC_12_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_25, data_out=>output_MAC_12_25);

	MAC_12_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_26, data_out=>output_MAC_12_26);

	MAC_12_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_27, data_out=>output_MAC_12_27);

	MAC_12_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_28, data_out=>output_MAC_12_28);

	MAC_12_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_29, data_out=>output_MAC_12_29);

	MAC_12_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_30, data_out=>output_MAC_12_30);

	MAC_12_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_12, data_in_B=>reg_input_col_31, data_out=>output_MAC_12_31);

	MAC_13_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_0, data_out=>output_MAC_13_0);

	MAC_13_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_1, data_out=>output_MAC_13_1);

	MAC_13_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_2, data_out=>output_MAC_13_2);

	MAC_13_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_3, data_out=>output_MAC_13_3);

	MAC_13_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_4, data_out=>output_MAC_13_4);

	MAC_13_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_5, data_out=>output_MAC_13_5);

	MAC_13_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_6, data_out=>output_MAC_13_6);

	MAC_13_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_7, data_out=>output_MAC_13_7);

	MAC_13_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_8, data_out=>output_MAC_13_8);

	MAC_13_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_9, data_out=>output_MAC_13_9);

	MAC_13_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_10, data_out=>output_MAC_13_10);

	MAC_13_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_11, data_out=>output_MAC_13_11);

	MAC_13_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_12, data_out=>output_MAC_13_12);

	MAC_13_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_13, data_out=>output_MAC_13_13);

	MAC_13_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_14, data_out=>output_MAC_13_14);

	MAC_13_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_15, data_out=>output_MAC_13_15);

	MAC_13_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_16, data_out=>output_MAC_13_16);

	MAC_13_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_17, data_out=>output_MAC_13_17);

	MAC_13_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_18, data_out=>output_MAC_13_18);

	MAC_13_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_19, data_out=>output_MAC_13_19);

	MAC_13_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_20, data_out=>output_MAC_13_20);

	MAC_13_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_21, data_out=>output_MAC_13_21);

	MAC_13_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_22, data_out=>output_MAC_13_22);

	MAC_13_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_23, data_out=>output_MAC_13_23);

	MAC_13_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_24, data_out=>output_MAC_13_24);

	MAC_13_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_25, data_out=>output_MAC_13_25);

	MAC_13_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_26, data_out=>output_MAC_13_26);

	MAC_13_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_27, data_out=>output_MAC_13_27);

	MAC_13_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_28, data_out=>output_MAC_13_28);

	MAC_13_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_29, data_out=>output_MAC_13_29);

	MAC_13_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_30, data_out=>output_MAC_13_30);

	MAC_13_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_13, data_in_B=>reg_input_col_31, data_out=>output_MAC_13_31);

	MAC_14_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_0, data_out=>output_MAC_14_0);

	MAC_14_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_1, data_out=>output_MAC_14_1);

	MAC_14_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_2, data_out=>output_MAC_14_2);

	MAC_14_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_3, data_out=>output_MAC_14_3);

	MAC_14_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_4, data_out=>output_MAC_14_4);

	MAC_14_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_5, data_out=>output_MAC_14_5);

	MAC_14_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_6, data_out=>output_MAC_14_6);

	MAC_14_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_7, data_out=>output_MAC_14_7);

	MAC_14_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_8, data_out=>output_MAC_14_8);

	MAC_14_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_9, data_out=>output_MAC_14_9);

	MAC_14_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_10, data_out=>output_MAC_14_10);

	MAC_14_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_11, data_out=>output_MAC_14_11);

	MAC_14_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_12, data_out=>output_MAC_14_12);

	MAC_14_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_13, data_out=>output_MAC_14_13);

	MAC_14_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_14, data_out=>output_MAC_14_14);

	MAC_14_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_15, data_out=>output_MAC_14_15);

	MAC_14_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_16, data_out=>output_MAC_14_16);

	MAC_14_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_17, data_out=>output_MAC_14_17);

	MAC_14_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_18, data_out=>output_MAC_14_18);

	MAC_14_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_19, data_out=>output_MAC_14_19);

	MAC_14_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_20, data_out=>output_MAC_14_20);

	MAC_14_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_21, data_out=>output_MAC_14_21);

	MAC_14_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_22, data_out=>output_MAC_14_22);

	MAC_14_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_23, data_out=>output_MAC_14_23);

	MAC_14_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_24, data_out=>output_MAC_14_24);

	MAC_14_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_25, data_out=>output_MAC_14_25);

	MAC_14_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_26, data_out=>output_MAC_14_26);

	MAC_14_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_27, data_out=>output_MAC_14_27);

	MAC_14_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_28, data_out=>output_MAC_14_28);

	MAC_14_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_29, data_out=>output_MAC_14_29);

	MAC_14_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_30, data_out=>output_MAC_14_30);

	MAC_14_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_14, data_in_B=>reg_input_col_31, data_out=>output_MAC_14_31);

	MAC_15_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_0, data_out=>output_MAC_15_0);

	MAC_15_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_1, data_out=>output_MAC_15_1);

	MAC_15_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_2, data_out=>output_MAC_15_2);

	MAC_15_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_3, data_out=>output_MAC_15_3);

	MAC_15_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_4, data_out=>output_MAC_15_4);

	MAC_15_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_5, data_out=>output_MAC_15_5);

	MAC_15_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_6, data_out=>output_MAC_15_6);

	MAC_15_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_7, data_out=>output_MAC_15_7);

	MAC_15_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_8, data_out=>output_MAC_15_8);

	MAC_15_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_9, data_out=>output_MAC_15_9);

	MAC_15_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_10, data_out=>output_MAC_15_10);

	MAC_15_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_11, data_out=>output_MAC_15_11);

	MAC_15_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_12, data_out=>output_MAC_15_12);

	MAC_15_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_13, data_out=>output_MAC_15_13);

	MAC_15_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_14, data_out=>output_MAC_15_14);

	MAC_15_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_15, data_out=>output_MAC_15_15);

	MAC_15_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_16, data_out=>output_MAC_15_16);

	MAC_15_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_17, data_out=>output_MAC_15_17);

	MAC_15_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_18, data_out=>output_MAC_15_18);

	MAC_15_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_19, data_out=>output_MAC_15_19);

	MAC_15_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_20, data_out=>output_MAC_15_20);

	MAC_15_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_21, data_out=>output_MAC_15_21);

	MAC_15_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_22, data_out=>output_MAC_15_22);

	MAC_15_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_23, data_out=>output_MAC_15_23);

	MAC_15_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_24, data_out=>output_MAC_15_24);

	MAC_15_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_25, data_out=>output_MAC_15_25);

	MAC_15_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_26, data_out=>output_MAC_15_26);

	MAC_15_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_27, data_out=>output_MAC_15_27);

	MAC_15_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_28, data_out=>output_MAC_15_28);

	MAC_15_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_29, data_out=>output_MAC_15_29);

	MAC_15_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_30, data_out=>output_MAC_15_30);

	MAC_15_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_15, data_in_B=>reg_input_col_31, data_out=>output_MAC_15_31);

	MAC_16_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_0, data_out=>output_MAC_16_0);

	MAC_16_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_1, data_out=>output_MAC_16_1);

	MAC_16_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_2, data_out=>output_MAC_16_2);

	MAC_16_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_3, data_out=>output_MAC_16_3);

	MAC_16_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_4, data_out=>output_MAC_16_4);

	MAC_16_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_5, data_out=>output_MAC_16_5);

	MAC_16_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_6, data_out=>output_MAC_16_6);

	MAC_16_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_7, data_out=>output_MAC_16_7);

	MAC_16_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_8, data_out=>output_MAC_16_8);

	MAC_16_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_9, data_out=>output_MAC_16_9);

	MAC_16_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_10, data_out=>output_MAC_16_10);

	MAC_16_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_11, data_out=>output_MAC_16_11);

	MAC_16_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_12, data_out=>output_MAC_16_12);

	MAC_16_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_13, data_out=>output_MAC_16_13);

	MAC_16_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_14, data_out=>output_MAC_16_14);

	MAC_16_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_15, data_out=>output_MAC_16_15);

	MAC_16_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_16, data_out=>output_MAC_16_16);

	MAC_16_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_17, data_out=>output_MAC_16_17);

	MAC_16_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_18, data_out=>output_MAC_16_18);

	MAC_16_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_19, data_out=>output_MAC_16_19);

	MAC_16_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_20, data_out=>output_MAC_16_20);

	MAC_16_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_21, data_out=>output_MAC_16_21);

	MAC_16_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_22, data_out=>output_MAC_16_22);

	MAC_16_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_23, data_out=>output_MAC_16_23);

	MAC_16_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_24, data_out=>output_MAC_16_24);

	MAC_16_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_25, data_out=>output_MAC_16_25);

	MAC_16_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_26, data_out=>output_MAC_16_26);

	MAC_16_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_27, data_out=>output_MAC_16_27);

	MAC_16_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_28, data_out=>output_MAC_16_28);

	MAC_16_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_29, data_out=>output_MAC_16_29);

	MAC_16_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_30, data_out=>output_MAC_16_30);

	MAC_16_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_16, data_in_B=>reg_input_col_31, data_out=>output_MAC_16_31);

	MAC_17_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_0, data_out=>output_MAC_17_0);

	MAC_17_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_1, data_out=>output_MAC_17_1);

	MAC_17_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_2, data_out=>output_MAC_17_2);

	MAC_17_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_3, data_out=>output_MAC_17_3);

	MAC_17_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_4, data_out=>output_MAC_17_4);

	MAC_17_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_5, data_out=>output_MAC_17_5);

	MAC_17_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_6, data_out=>output_MAC_17_6);

	MAC_17_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_7, data_out=>output_MAC_17_7);

	MAC_17_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_8, data_out=>output_MAC_17_8);

	MAC_17_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_9, data_out=>output_MAC_17_9);

	MAC_17_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_10, data_out=>output_MAC_17_10);

	MAC_17_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_11, data_out=>output_MAC_17_11);

	MAC_17_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_12, data_out=>output_MAC_17_12);

	MAC_17_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_13, data_out=>output_MAC_17_13);

	MAC_17_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_14, data_out=>output_MAC_17_14);

	MAC_17_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_15, data_out=>output_MAC_17_15);

	MAC_17_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_16, data_out=>output_MAC_17_16);

	MAC_17_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_17, data_out=>output_MAC_17_17);

	MAC_17_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_18, data_out=>output_MAC_17_18);

	MAC_17_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_19, data_out=>output_MAC_17_19);

	MAC_17_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_20, data_out=>output_MAC_17_20);

	MAC_17_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_21, data_out=>output_MAC_17_21);

	MAC_17_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_22, data_out=>output_MAC_17_22);

	MAC_17_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_23, data_out=>output_MAC_17_23);

	MAC_17_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_24, data_out=>output_MAC_17_24);

	MAC_17_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_25, data_out=>output_MAC_17_25);

	MAC_17_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_26, data_out=>output_MAC_17_26);

	MAC_17_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_27, data_out=>output_MAC_17_27);

	MAC_17_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_28, data_out=>output_MAC_17_28);

	MAC_17_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_29, data_out=>output_MAC_17_29);

	MAC_17_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_30, data_out=>output_MAC_17_30);

	MAC_17_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_17, data_in_B=>reg_input_col_31, data_out=>output_MAC_17_31);

	MAC_18_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_0, data_out=>output_MAC_18_0);

	MAC_18_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_1, data_out=>output_MAC_18_1);

	MAC_18_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_2, data_out=>output_MAC_18_2);

	MAC_18_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_3, data_out=>output_MAC_18_3);

	MAC_18_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_4, data_out=>output_MAC_18_4);

	MAC_18_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_5, data_out=>output_MAC_18_5);

	MAC_18_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_6, data_out=>output_MAC_18_6);

	MAC_18_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_7, data_out=>output_MAC_18_7);

	MAC_18_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_8, data_out=>output_MAC_18_8);

	MAC_18_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_9, data_out=>output_MAC_18_9);

	MAC_18_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_10, data_out=>output_MAC_18_10);

	MAC_18_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_11, data_out=>output_MAC_18_11);

	MAC_18_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_12, data_out=>output_MAC_18_12);

	MAC_18_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_13, data_out=>output_MAC_18_13);

	MAC_18_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_14, data_out=>output_MAC_18_14);

	MAC_18_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_15, data_out=>output_MAC_18_15);

	MAC_18_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_16, data_out=>output_MAC_18_16);

	MAC_18_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_17, data_out=>output_MAC_18_17);

	MAC_18_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_18, data_out=>output_MAC_18_18);

	MAC_18_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_19, data_out=>output_MAC_18_19);

	MAC_18_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_20, data_out=>output_MAC_18_20);

	MAC_18_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_21, data_out=>output_MAC_18_21);

	MAC_18_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_22, data_out=>output_MAC_18_22);

	MAC_18_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_23, data_out=>output_MAC_18_23);

	MAC_18_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_24, data_out=>output_MAC_18_24);

	MAC_18_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_25, data_out=>output_MAC_18_25);

	MAC_18_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_26, data_out=>output_MAC_18_26);

	MAC_18_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_27, data_out=>output_MAC_18_27);

	MAC_18_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_28, data_out=>output_MAC_18_28);

	MAC_18_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_29, data_out=>output_MAC_18_29);

	MAC_18_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_30, data_out=>output_MAC_18_30);

	MAC_18_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_18, data_in_B=>reg_input_col_31, data_out=>output_MAC_18_31);

	MAC_19_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_0, data_out=>output_MAC_19_0);

	MAC_19_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_1, data_out=>output_MAC_19_1);

	MAC_19_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_2, data_out=>output_MAC_19_2);

	MAC_19_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_3, data_out=>output_MAC_19_3);

	MAC_19_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_4, data_out=>output_MAC_19_4);

	MAC_19_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_5, data_out=>output_MAC_19_5);

	MAC_19_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_6, data_out=>output_MAC_19_6);

	MAC_19_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_7, data_out=>output_MAC_19_7);

	MAC_19_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_8, data_out=>output_MAC_19_8);

	MAC_19_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_9, data_out=>output_MAC_19_9);

	MAC_19_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_10, data_out=>output_MAC_19_10);

	MAC_19_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_11, data_out=>output_MAC_19_11);

	MAC_19_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_12, data_out=>output_MAC_19_12);

	MAC_19_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_13, data_out=>output_MAC_19_13);

	MAC_19_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_14, data_out=>output_MAC_19_14);

	MAC_19_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_15, data_out=>output_MAC_19_15);

	MAC_19_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_16, data_out=>output_MAC_19_16);

	MAC_19_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_17, data_out=>output_MAC_19_17);

	MAC_19_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_18, data_out=>output_MAC_19_18);

	MAC_19_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_19, data_out=>output_MAC_19_19);

	MAC_19_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_20, data_out=>output_MAC_19_20);

	MAC_19_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_21, data_out=>output_MAC_19_21);

	MAC_19_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_22, data_out=>output_MAC_19_22);

	MAC_19_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_23, data_out=>output_MAC_19_23);

	MAC_19_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_24, data_out=>output_MAC_19_24);

	MAC_19_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_25, data_out=>output_MAC_19_25);

	MAC_19_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_26, data_out=>output_MAC_19_26);

	MAC_19_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_27, data_out=>output_MAC_19_27);

	MAC_19_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_28, data_out=>output_MAC_19_28);

	MAC_19_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_29, data_out=>output_MAC_19_29);

	MAC_19_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_30, data_out=>output_MAC_19_30);

	MAC_19_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_19, data_in_B=>reg_input_col_31, data_out=>output_MAC_19_31);

	MAC_20_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_0, data_out=>output_MAC_20_0);

	MAC_20_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_1, data_out=>output_MAC_20_1);

	MAC_20_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_2, data_out=>output_MAC_20_2);

	MAC_20_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_3, data_out=>output_MAC_20_3);

	MAC_20_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_4, data_out=>output_MAC_20_4);

	MAC_20_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_5, data_out=>output_MAC_20_5);

	MAC_20_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_6, data_out=>output_MAC_20_6);

	MAC_20_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_7, data_out=>output_MAC_20_7);

	MAC_20_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_8, data_out=>output_MAC_20_8);

	MAC_20_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_9, data_out=>output_MAC_20_9);

	MAC_20_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_10, data_out=>output_MAC_20_10);

	MAC_20_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_11, data_out=>output_MAC_20_11);

	MAC_20_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_12, data_out=>output_MAC_20_12);

	MAC_20_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_13, data_out=>output_MAC_20_13);

	MAC_20_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_14, data_out=>output_MAC_20_14);

	MAC_20_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_15, data_out=>output_MAC_20_15);

	MAC_20_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_16, data_out=>output_MAC_20_16);

	MAC_20_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_17, data_out=>output_MAC_20_17);

	MAC_20_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_18, data_out=>output_MAC_20_18);

	MAC_20_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_19, data_out=>output_MAC_20_19);

	MAC_20_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_20, data_out=>output_MAC_20_20);

	MAC_20_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_21, data_out=>output_MAC_20_21);

	MAC_20_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_22, data_out=>output_MAC_20_22);

	MAC_20_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_23, data_out=>output_MAC_20_23);

	MAC_20_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_24, data_out=>output_MAC_20_24);

	MAC_20_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_25, data_out=>output_MAC_20_25);

	MAC_20_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_26, data_out=>output_MAC_20_26);

	MAC_20_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_27, data_out=>output_MAC_20_27);

	MAC_20_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_28, data_out=>output_MAC_20_28);

	MAC_20_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_29, data_out=>output_MAC_20_29);

	MAC_20_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_30, data_out=>output_MAC_20_30);

	MAC_20_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_20, data_in_B=>reg_input_col_31, data_out=>output_MAC_20_31);

	MAC_21_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_0, data_out=>output_MAC_21_0);

	MAC_21_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_1, data_out=>output_MAC_21_1);

	MAC_21_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_2, data_out=>output_MAC_21_2);

	MAC_21_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_3, data_out=>output_MAC_21_3);

	MAC_21_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_4, data_out=>output_MAC_21_4);

	MAC_21_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_5, data_out=>output_MAC_21_5);

	MAC_21_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_6, data_out=>output_MAC_21_6);

	MAC_21_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_7, data_out=>output_MAC_21_7);

	MAC_21_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_8, data_out=>output_MAC_21_8);

	MAC_21_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_9, data_out=>output_MAC_21_9);

	MAC_21_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_10, data_out=>output_MAC_21_10);

	MAC_21_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_11, data_out=>output_MAC_21_11);

	MAC_21_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_12, data_out=>output_MAC_21_12);

	MAC_21_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_13, data_out=>output_MAC_21_13);

	MAC_21_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_14, data_out=>output_MAC_21_14);

	MAC_21_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_15, data_out=>output_MAC_21_15);

	MAC_21_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_16, data_out=>output_MAC_21_16);

	MAC_21_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_17, data_out=>output_MAC_21_17);

	MAC_21_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_18, data_out=>output_MAC_21_18);

	MAC_21_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_19, data_out=>output_MAC_21_19);

	MAC_21_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_20, data_out=>output_MAC_21_20);

	MAC_21_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_21, data_out=>output_MAC_21_21);

	MAC_21_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_22, data_out=>output_MAC_21_22);

	MAC_21_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_23, data_out=>output_MAC_21_23);

	MAC_21_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_24, data_out=>output_MAC_21_24);

	MAC_21_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_25, data_out=>output_MAC_21_25);

	MAC_21_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_26, data_out=>output_MAC_21_26);

	MAC_21_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_27, data_out=>output_MAC_21_27);

	MAC_21_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_28, data_out=>output_MAC_21_28);

	MAC_21_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_29, data_out=>output_MAC_21_29);

	MAC_21_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_30, data_out=>output_MAC_21_30);

	MAC_21_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_21, data_in_B=>reg_input_col_31, data_out=>output_MAC_21_31);

	MAC_22_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_0, data_out=>output_MAC_22_0);

	MAC_22_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_1, data_out=>output_MAC_22_1);

	MAC_22_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_2, data_out=>output_MAC_22_2);

	MAC_22_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_3, data_out=>output_MAC_22_3);

	MAC_22_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_4, data_out=>output_MAC_22_4);

	MAC_22_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_5, data_out=>output_MAC_22_5);

	MAC_22_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_6, data_out=>output_MAC_22_6);

	MAC_22_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_7, data_out=>output_MAC_22_7);

	MAC_22_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_8, data_out=>output_MAC_22_8);

	MAC_22_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_9, data_out=>output_MAC_22_9);

	MAC_22_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_10, data_out=>output_MAC_22_10);

	MAC_22_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_11, data_out=>output_MAC_22_11);

	MAC_22_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_12, data_out=>output_MAC_22_12);

	MAC_22_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_13, data_out=>output_MAC_22_13);

	MAC_22_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_14, data_out=>output_MAC_22_14);

	MAC_22_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_15, data_out=>output_MAC_22_15);

	MAC_22_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_16, data_out=>output_MAC_22_16);

	MAC_22_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_17, data_out=>output_MAC_22_17);

	MAC_22_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_18, data_out=>output_MAC_22_18);

	MAC_22_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_19, data_out=>output_MAC_22_19);

	MAC_22_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_20, data_out=>output_MAC_22_20);

	MAC_22_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_21, data_out=>output_MAC_22_21);

	MAC_22_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_22, data_out=>output_MAC_22_22);

	MAC_22_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_23, data_out=>output_MAC_22_23);

	MAC_22_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_24, data_out=>output_MAC_22_24);

	MAC_22_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_25, data_out=>output_MAC_22_25);

	MAC_22_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_26, data_out=>output_MAC_22_26);

	MAC_22_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_27, data_out=>output_MAC_22_27);

	MAC_22_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_28, data_out=>output_MAC_22_28);

	MAC_22_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_29, data_out=>output_MAC_22_29);

	MAC_22_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_30, data_out=>output_MAC_22_30);

	MAC_22_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_22, data_in_B=>reg_input_col_31, data_out=>output_MAC_22_31);

	MAC_23_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_0, data_out=>output_MAC_23_0);

	MAC_23_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_1, data_out=>output_MAC_23_1);

	MAC_23_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_2, data_out=>output_MAC_23_2);

	MAC_23_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_3, data_out=>output_MAC_23_3);

	MAC_23_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_4, data_out=>output_MAC_23_4);

	MAC_23_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_5, data_out=>output_MAC_23_5);

	MAC_23_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_6, data_out=>output_MAC_23_6);

	MAC_23_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_7, data_out=>output_MAC_23_7);

	MAC_23_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_8, data_out=>output_MAC_23_8);

	MAC_23_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_9, data_out=>output_MAC_23_9);

	MAC_23_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_10, data_out=>output_MAC_23_10);

	MAC_23_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_11, data_out=>output_MAC_23_11);

	MAC_23_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_12, data_out=>output_MAC_23_12);

	MAC_23_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_13, data_out=>output_MAC_23_13);

	MAC_23_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_14, data_out=>output_MAC_23_14);

	MAC_23_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_15, data_out=>output_MAC_23_15);

	MAC_23_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_16, data_out=>output_MAC_23_16);

	MAC_23_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_17, data_out=>output_MAC_23_17);

	MAC_23_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_18, data_out=>output_MAC_23_18);

	MAC_23_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_19, data_out=>output_MAC_23_19);

	MAC_23_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_20, data_out=>output_MAC_23_20);

	MAC_23_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_21, data_out=>output_MAC_23_21);

	MAC_23_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_22, data_out=>output_MAC_23_22);

	MAC_23_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_23, data_out=>output_MAC_23_23);

	MAC_23_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_24, data_out=>output_MAC_23_24);

	MAC_23_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_25, data_out=>output_MAC_23_25);

	MAC_23_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_26, data_out=>output_MAC_23_26);

	MAC_23_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_27, data_out=>output_MAC_23_27);

	MAC_23_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_28, data_out=>output_MAC_23_28);

	MAC_23_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_29, data_out=>output_MAC_23_29);

	MAC_23_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_30, data_out=>output_MAC_23_30);

	MAC_23_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_23, data_in_B=>reg_input_col_31, data_out=>output_MAC_23_31);

	MAC_24_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_0, data_out=>output_MAC_24_0);

	MAC_24_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_1, data_out=>output_MAC_24_1);

	MAC_24_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_2, data_out=>output_MAC_24_2);

	MAC_24_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_3, data_out=>output_MAC_24_3);

	MAC_24_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_4, data_out=>output_MAC_24_4);

	MAC_24_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_5, data_out=>output_MAC_24_5);

	MAC_24_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_6, data_out=>output_MAC_24_6);

	MAC_24_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_7, data_out=>output_MAC_24_7);

	MAC_24_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_8, data_out=>output_MAC_24_8);

	MAC_24_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_9, data_out=>output_MAC_24_9);

	MAC_24_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_10, data_out=>output_MAC_24_10);

	MAC_24_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_11, data_out=>output_MAC_24_11);

	MAC_24_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_12, data_out=>output_MAC_24_12);

	MAC_24_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_13, data_out=>output_MAC_24_13);

	MAC_24_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_14, data_out=>output_MAC_24_14);

	MAC_24_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_15, data_out=>output_MAC_24_15);

	MAC_24_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_16, data_out=>output_MAC_24_16);

	MAC_24_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_17, data_out=>output_MAC_24_17);

	MAC_24_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_18, data_out=>output_MAC_24_18);

	MAC_24_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_19, data_out=>output_MAC_24_19);

	MAC_24_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_20, data_out=>output_MAC_24_20);

	MAC_24_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_21, data_out=>output_MAC_24_21);

	MAC_24_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_22, data_out=>output_MAC_24_22);

	MAC_24_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_23, data_out=>output_MAC_24_23);

	MAC_24_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_24, data_out=>output_MAC_24_24);

	MAC_24_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_25, data_out=>output_MAC_24_25);

	MAC_24_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_26, data_out=>output_MAC_24_26);

	MAC_24_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_27, data_out=>output_MAC_24_27);

	MAC_24_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_28, data_out=>output_MAC_24_28);

	MAC_24_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_29, data_out=>output_MAC_24_29);

	MAC_24_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_30, data_out=>output_MAC_24_30);

	MAC_24_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_24, data_in_B=>reg_input_col_31, data_out=>output_MAC_24_31);

	MAC_25_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_0, data_out=>output_MAC_25_0);

	MAC_25_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_1, data_out=>output_MAC_25_1);

	MAC_25_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_2, data_out=>output_MAC_25_2);

	MAC_25_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_3, data_out=>output_MAC_25_3);

	MAC_25_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_4, data_out=>output_MAC_25_4);

	MAC_25_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_5, data_out=>output_MAC_25_5);

	MAC_25_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_6, data_out=>output_MAC_25_6);

	MAC_25_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_7, data_out=>output_MAC_25_7);

	MAC_25_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_8, data_out=>output_MAC_25_8);

	MAC_25_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_9, data_out=>output_MAC_25_9);

	MAC_25_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_10, data_out=>output_MAC_25_10);

	MAC_25_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_11, data_out=>output_MAC_25_11);

	MAC_25_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_12, data_out=>output_MAC_25_12);

	MAC_25_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_13, data_out=>output_MAC_25_13);

	MAC_25_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_14, data_out=>output_MAC_25_14);

	MAC_25_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_15, data_out=>output_MAC_25_15);

	MAC_25_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_16, data_out=>output_MAC_25_16);

	MAC_25_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_17, data_out=>output_MAC_25_17);

	MAC_25_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_18, data_out=>output_MAC_25_18);

	MAC_25_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_19, data_out=>output_MAC_25_19);

	MAC_25_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_20, data_out=>output_MAC_25_20);

	MAC_25_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_21, data_out=>output_MAC_25_21);

	MAC_25_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_22, data_out=>output_MAC_25_22);

	MAC_25_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_23, data_out=>output_MAC_25_23);

	MAC_25_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_24, data_out=>output_MAC_25_24);

	MAC_25_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_25, data_out=>output_MAC_25_25);

	MAC_25_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_26, data_out=>output_MAC_25_26);

	MAC_25_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_27, data_out=>output_MAC_25_27);

	MAC_25_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_28, data_out=>output_MAC_25_28);

	MAC_25_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_29, data_out=>output_MAC_25_29);

	MAC_25_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_30, data_out=>output_MAC_25_30);

	MAC_25_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_25, data_in_B=>reg_input_col_31, data_out=>output_MAC_25_31);

	MAC_26_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_0, data_out=>output_MAC_26_0);

	MAC_26_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_1, data_out=>output_MAC_26_1);

	MAC_26_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_2, data_out=>output_MAC_26_2);

	MAC_26_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_3, data_out=>output_MAC_26_3);

	MAC_26_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_4, data_out=>output_MAC_26_4);

	MAC_26_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_5, data_out=>output_MAC_26_5);

	MAC_26_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_6, data_out=>output_MAC_26_6);

	MAC_26_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_7, data_out=>output_MAC_26_7);

	MAC_26_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_8, data_out=>output_MAC_26_8);

	MAC_26_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_9, data_out=>output_MAC_26_9);

	MAC_26_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_10, data_out=>output_MAC_26_10);

	MAC_26_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_11, data_out=>output_MAC_26_11);

	MAC_26_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_12, data_out=>output_MAC_26_12);

	MAC_26_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_13, data_out=>output_MAC_26_13);

	MAC_26_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_14, data_out=>output_MAC_26_14);

	MAC_26_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_15, data_out=>output_MAC_26_15);

	MAC_26_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_16, data_out=>output_MAC_26_16);

	MAC_26_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_17, data_out=>output_MAC_26_17);

	MAC_26_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_18, data_out=>output_MAC_26_18);

	MAC_26_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_19, data_out=>output_MAC_26_19);

	MAC_26_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_20, data_out=>output_MAC_26_20);

	MAC_26_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_21, data_out=>output_MAC_26_21);

	MAC_26_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_22, data_out=>output_MAC_26_22);

	MAC_26_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_23, data_out=>output_MAC_26_23);

	MAC_26_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_24, data_out=>output_MAC_26_24);

	MAC_26_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_25, data_out=>output_MAC_26_25);

	MAC_26_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_26, data_out=>output_MAC_26_26);

	MAC_26_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_27, data_out=>output_MAC_26_27);

	MAC_26_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_28, data_out=>output_MAC_26_28);

	MAC_26_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_29, data_out=>output_MAC_26_29);

	MAC_26_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_30, data_out=>output_MAC_26_30);

	MAC_26_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_26, data_in_B=>reg_input_col_31, data_out=>output_MAC_26_31);

	MAC_27_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_0, data_out=>output_MAC_27_0);

	MAC_27_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_1, data_out=>output_MAC_27_1);

	MAC_27_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_2, data_out=>output_MAC_27_2);

	MAC_27_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_3, data_out=>output_MAC_27_3);

	MAC_27_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_4, data_out=>output_MAC_27_4);

	MAC_27_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_5, data_out=>output_MAC_27_5);

	MAC_27_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_6, data_out=>output_MAC_27_6);

	MAC_27_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_7, data_out=>output_MAC_27_7);

	MAC_27_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_8, data_out=>output_MAC_27_8);

	MAC_27_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_9, data_out=>output_MAC_27_9);

	MAC_27_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_10, data_out=>output_MAC_27_10);

	MAC_27_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_11, data_out=>output_MAC_27_11);

	MAC_27_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_12, data_out=>output_MAC_27_12);

	MAC_27_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_13, data_out=>output_MAC_27_13);

	MAC_27_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_14, data_out=>output_MAC_27_14);

	MAC_27_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_15, data_out=>output_MAC_27_15);

	MAC_27_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_16, data_out=>output_MAC_27_16);

	MAC_27_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_17, data_out=>output_MAC_27_17);

	MAC_27_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_18, data_out=>output_MAC_27_18);

	MAC_27_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_19, data_out=>output_MAC_27_19);

	MAC_27_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_20, data_out=>output_MAC_27_20);

	MAC_27_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_21, data_out=>output_MAC_27_21);

	MAC_27_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_22, data_out=>output_MAC_27_22);

	MAC_27_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_23, data_out=>output_MAC_27_23);

	MAC_27_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_24, data_out=>output_MAC_27_24);

	MAC_27_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_25, data_out=>output_MAC_27_25);

	MAC_27_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_26, data_out=>output_MAC_27_26);

	MAC_27_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_27, data_out=>output_MAC_27_27);

	MAC_27_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_28, data_out=>output_MAC_27_28);

	MAC_27_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_29, data_out=>output_MAC_27_29);

	MAC_27_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_30, data_out=>output_MAC_27_30);

	MAC_27_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_27, data_in_B=>reg_input_col_31, data_out=>output_MAC_27_31);

	MAC_28_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_0, data_out=>output_MAC_28_0);

	MAC_28_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_1, data_out=>output_MAC_28_1);

	MAC_28_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_2, data_out=>output_MAC_28_2);

	MAC_28_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_3, data_out=>output_MAC_28_3);

	MAC_28_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_4, data_out=>output_MAC_28_4);

	MAC_28_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_5, data_out=>output_MAC_28_5);

	MAC_28_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_6, data_out=>output_MAC_28_6);

	MAC_28_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_7, data_out=>output_MAC_28_7);

	MAC_28_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_8, data_out=>output_MAC_28_8);

	MAC_28_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_9, data_out=>output_MAC_28_9);

	MAC_28_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_10, data_out=>output_MAC_28_10);

	MAC_28_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_11, data_out=>output_MAC_28_11);

	MAC_28_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_12, data_out=>output_MAC_28_12);

	MAC_28_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_13, data_out=>output_MAC_28_13);

	MAC_28_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_14, data_out=>output_MAC_28_14);

	MAC_28_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_15, data_out=>output_MAC_28_15);

	MAC_28_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_16, data_out=>output_MAC_28_16);

	MAC_28_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_17, data_out=>output_MAC_28_17);

	MAC_28_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_18, data_out=>output_MAC_28_18);

	MAC_28_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_19, data_out=>output_MAC_28_19);

	MAC_28_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_20, data_out=>output_MAC_28_20);

	MAC_28_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_21, data_out=>output_MAC_28_21);

	MAC_28_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_22, data_out=>output_MAC_28_22);

	MAC_28_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_23, data_out=>output_MAC_28_23);

	MAC_28_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_24, data_out=>output_MAC_28_24);

	MAC_28_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_25, data_out=>output_MAC_28_25);

	MAC_28_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_26, data_out=>output_MAC_28_26);

	MAC_28_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_27, data_out=>output_MAC_28_27);

	MAC_28_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_28, data_out=>output_MAC_28_28);

	MAC_28_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_29, data_out=>output_MAC_28_29);

	MAC_28_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_30, data_out=>output_MAC_28_30);

	MAC_28_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_28, data_in_B=>reg_input_col_31, data_out=>output_MAC_28_31);

	MAC_29_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_0, data_out=>output_MAC_29_0);

	MAC_29_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_1, data_out=>output_MAC_29_1);

	MAC_29_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_2, data_out=>output_MAC_29_2);

	MAC_29_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_3, data_out=>output_MAC_29_3);

	MAC_29_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_4, data_out=>output_MAC_29_4);

	MAC_29_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_5, data_out=>output_MAC_29_5);

	MAC_29_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_6, data_out=>output_MAC_29_6);

	MAC_29_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_7, data_out=>output_MAC_29_7);

	MAC_29_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_8, data_out=>output_MAC_29_8);

	MAC_29_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_9, data_out=>output_MAC_29_9);

	MAC_29_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_10, data_out=>output_MAC_29_10);

	MAC_29_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_11, data_out=>output_MAC_29_11);

	MAC_29_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_12, data_out=>output_MAC_29_12);

	MAC_29_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_13, data_out=>output_MAC_29_13);

	MAC_29_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_14, data_out=>output_MAC_29_14);

	MAC_29_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_15, data_out=>output_MAC_29_15);

	MAC_29_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_16, data_out=>output_MAC_29_16);

	MAC_29_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_17, data_out=>output_MAC_29_17);

	MAC_29_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_18, data_out=>output_MAC_29_18);

	MAC_29_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_19, data_out=>output_MAC_29_19);

	MAC_29_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_20, data_out=>output_MAC_29_20);

	MAC_29_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_21, data_out=>output_MAC_29_21);

	MAC_29_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_22, data_out=>output_MAC_29_22);

	MAC_29_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_23, data_out=>output_MAC_29_23);

	MAC_29_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_24, data_out=>output_MAC_29_24);

	MAC_29_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_25, data_out=>output_MAC_29_25);

	MAC_29_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_26, data_out=>output_MAC_29_26);

	MAC_29_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_27, data_out=>output_MAC_29_27);

	MAC_29_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_28, data_out=>output_MAC_29_28);

	MAC_29_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_29, data_out=>output_MAC_29_29);

	MAC_29_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_30, data_out=>output_MAC_29_30);

	MAC_29_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_29, data_in_B=>reg_input_col_31, data_out=>output_MAC_29_31);

	MAC_30_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_0, data_out=>output_MAC_30_0);

	MAC_30_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_1, data_out=>output_MAC_30_1);

	MAC_30_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_2, data_out=>output_MAC_30_2);

	MAC_30_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_3, data_out=>output_MAC_30_3);

	MAC_30_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_4, data_out=>output_MAC_30_4);

	MAC_30_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_5, data_out=>output_MAC_30_5);

	MAC_30_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_6, data_out=>output_MAC_30_6);

	MAC_30_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_7, data_out=>output_MAC_30_7);

	MAC_30_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_8, data_out=>output_MAC_30_8);

	MAC_30_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_9, data_out=>output_MAC_30_9);

	MAC_30_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_10, data_out=>output_MAC_30_10);

	MAC_30_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_11, data_out=>output_MAC_30_11);

	MAC_30_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_12, data_out=>output_MAC_30_12);

	MAC_30_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_13, data_out=>output_MAC_30_13);

	MAC_30_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_14, data_out=>output_MAC_30_14);

	MAC_30_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_15, data_out=>output_MAC_30_15);

	MAC_30_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_16, data_out=>output_MAC_30_16);

	MAC_30_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_17, data_out=>output_MAC_30_17);

	MAC_30_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_18, data_out=>output_MAC_30_18);

	MAC_30_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_19, data_out=>output_MAC_30_19);

	MAC_30_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_20, data_out=>output_MAC_30_20);

	MAC_30_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_21, data_out=>output_MAC_30_21);

	MAC_30_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_22, data_out=>output_MAC_30_22);

	MAC_30_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_23, data_out=>output_MAC_30_23);

	MAC_30_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_24, data_out=>output_MAC_30_24);

	MAC_30_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_25, data_out=>output_MAC_30_25);

	MAC_30_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_26, data_out=>output_MAC_30_26);

	MAC_30_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_27, data_out=>output_MAC_30_27);

	MAC_30_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_28, data_out=>output_MAC_30_28);

	MAC_30_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_29, data_out=>output_MAC_30_29);

	MAC_30_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_30, data_out=>output_MAC_30_30);

	MAC_30_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_30, data_in_B=>reg_input_col_31, data_out=>output_MAC_30_31);

	MAC_31_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_0, data_out=>output_MAC_31_0);

	MAC_31_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_1, data_out=>output_MAC_31_1);

	MAC_31_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_2, data_out=>output_MAC_31_2);

	MAC_31_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_3, data_out=>output_MAC_31_3);

	MAC_31_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_4, data_out=>output_MAC_31_4);

	MAC_31_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_5, data_out=>output_MAC_31_5);

	MAC_31_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_6, data_out=>output_MAC_31_6);

	MAC_31_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_7, data_out=>output_MAC_31_7);

	MAC_31_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_8, data_out=>output_MAC_31_8);

	MAC_31_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_9, data_out=>output_MAC_31_9);

	MAC_31_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_10, data_out=>output_MAC_31_10);

	MAC_31_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_11, data_out=>output_MAC_31_11);

	MAC_31_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_12, data_out=>output_MAC_31_12);

	MAC_31_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_13, data_out=>output_MAC_31_13);

	MAC_31_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_14, data_out=>output_MAC_31_14);

	MAC_31_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_15, data_out=>output_MAC_31_15);

	MAC_31_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_16, data_out=>output_MAC_31_16);

	MAC_31_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_17, data_out=>output_MAC_31_17);

	MAC_31_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_18, data_out=>output_MAC_31_18);

	MAC_31_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_19, data_out=>output_MAC_31_19);

	MAC_31_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_20, data_out=>output_MAC_31_20);

	MAC_31_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_21, data_out=>output_MAC_31_21);

	MAC_31_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_22, data_out=>output_MAC_31_22);

	MAC_31_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_23, data_out=>output_MAC_31_23);

	MAC_31_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_24, data_out=>output_MAC_31_24);

	MAC_31_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_25, data_out=>output_MAC_31_25);

	MAC_31_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_26, data_out=>output_MAC_31_26);

	MAC_31_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_27, data_out=>output_MAC_31_27);

	MAC_31_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_28, data_out=>output_MAC_31_28);

	MAC_31_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_29, data_out=>output_MAC_31_29);

	MAC_31_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_30, data_out=>output_MAC_31_30);

	MAC_31_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>reg_ENABLE_in, data_in_A=>reg_input_row_31, data_in_B=>reg_input_col_31, data_out=>output_MAC_31_31);


	mux_row_0: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_0_0, I1=>output_MAC_0_1, I2=>output_MAC_0_2, I3=>output_MAC_0_3, I4=>output_MAC_0_4, I5=>output_MAC_0_5, I6=>output_MAC_0_6, I7=>output_MAC_0_7, I8=>output_MAC_0_8, I9=>output_MAC_0_9, I10=>output_MAC_0_10, I11=>output_MAC_0_11, I12=>output_MAC_0_12, I13=>output_MAC_0_13, I14=>output_MAC_0_14, I15=>output_MAC_0_15, I16=>output_MAC_0_16, I17=>output_MAC_0_17, I18=>output_MAC_0_18, I19=>output_MAC_0_19, I20=>output_MAC_0_20, I21=>output_MAC_0_21, I22=>output_MAC_0_22, I23=>output_MAC_0_23, I24=>output_MAC_0_24, I25=>output_MAC_0_25, I26=>output_MAC_0_26, I27=>output_MAC_0_27, I28=>output_MAC_0_28, I29=>output_MAC_0_29, I30=>output_MAC_0_30, I31=>output_MAC_0_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_0);

	mux_row_1: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_1_0, I1=>output_MAC_1_1, I2=>output_MAC_1_2, I3=>output_MAC_1_3, I4=>output_MAC_1_4, I5=>output_MAC_1_5, I6=>output_MAC_1_6, I7=>output_MAC_1_7, I8=>output_MAC_1_8, I9=>output_MAC_1_9, I10=>output_MAC_1_10, I11=>output_MAC_1_11, I12=>output_MAC_1_12, I13=>output_MAC_1_13, I14=>output_MAC_1_14, I15=>output_MAC_1_15, I16=>output_MAC_1_16, I17=>output_MAC_1_17, I18=>output_MAC_1_18, I19=>output_MAC_1_19, I20=>output_MAC_1_20, I21=>output_MAC_1_21, I22=>output_MAC_1_22, I23=>output_MAC_1_23, I24=>output_MAC_1_24, I25=>output_MAC_1_25, I26=>output_MAC_1_26, I27=>output_MAC_1_27, I28=>output_MAC_1_28, I29=>output_MAC_1_29, I30=>output_MAC_1_30, I31=>output_MAC_1_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_1);

	mux_row_2: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_2_0, I1=>output_MAC_2_1, I2=>output_MAC_2_2, I3=>output_MAC_2_3, I4=>output_MAC_2_4, I5=>output_MAC_2_5, I6=>output_MAC_2_6, I7=>output_MAC_2_7, I8=>output_MAC_2_8, I9=>output_MAC_2_9, I10=>output_MAC_2_10, I11=>output_MAC_2_11, I12=>output_MAC_2_12, I13=>output_MAC_2_13, I14=>output_MAC_2_14, I15=>output_MAC_2_15, I16=>output_MAC_2_16, I17=>output_MAC_2_17, I18=>output_MAC_2_18, I19=>output_MAC_2_19, I20=>output_MAC_2_20, I21=>output_MAC_2_21, I22=>output_MAC_2_22, I23=>output_MAC_2_23, I24=>output_MAC_2_24, I25=>output_MAC_2_25, I26=>output_MAC_2_26, I27=>output_MAC_2_27, I28=>output_MAC_2_28, I29=>output_MAC_2_29, I30=>output_MAC_2_30, I31=>output_MAC_2_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_2);

	mux_row_3: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_3_0, I1=>output_MAC_3_1, I2=>output_MAC_3_2, I3=>output_MAC_3_3, I4=>output_MAC_3_4, I5=>output_MAC_3_5, I6=>output_MAC_3_6, I7=>output_MAC_3_7, I8=>output_MAC_3_8, I9=>output_MAC_3_9, I10=>output_MAC_3_10, I11=>output_MAC_3_11, I12=>output_MAC_3_12, I13=>output_MAC_3_13, I14=>output_MAC_3_14, I15=>output_MAC_3_15, I16=>output_MAC_3_16, I17=>output_MAC_3_17, I18=>output_MAC_3_18, I19=>output_MAC_3_19, I20=>output_MAC_3_20, I21=>output_MAC_3_21, I22=>output_MAC_3_22, I23=>output_MAC_3_23, I24=>output_MAC_3_24, I25=>output_MAC_3_25, I26=>output_MAC_3_26, I27=>output_MAC_3_27, I28=>output_MAC_3_28, I29=>output_MAC_3_29, I30=>output_MAC_3_30, I31=>output_MAC_3_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_3);

	mux_row_4: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_4_0, I1=>output_MAC_4_1, I2=>output_MAC_4_2, I3=>output_MAC_4_3, I4=>output_MAC_4_4, I5=>output_MAC_4_5, I6=>output_MAC_4_6, I7=>output_MAC_4_7, I8=>output_MAC_4_8, I9=>output_MAC_4_9, I10=>output_MAC_4_10, I11=>output_MAC_4_11, I12=>output_MAC_4_12, I13=>output_MAC_4_13, I14=>output_MAC_4_14, I15=>output_MAC_4_15, I16=>output_MAC_4_16, I17=>output_MAC_4_17, I18=>output_MAC_4_18, I19=>output_MAC_4_19, I20=>output_MAC_4_20, I21=>output_MAC_4_21, I22=>output_MAC_4_22, I23=>output_MAC_4_23, I24=>output_MAC_4_24, I25=>output_MAC_4_25, I26=>output_MAC_4_26, I27=>output_MAC_4_27, I28=>output_MAC_4_28, I29=>output_MAC_4_29, I30=>output_MAC_4_30, I31=>output_MAC_4_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_4);

	mux_row_5: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_5_0, I1=>output_MAC_5_1, I2=>output_MAC_5_2, I3=>output_MAC_5_3, I4=>output_MAC_5_4, I5=>output_MAC_5_5, I6=>output_MAC_5_6, I7=>output_MAC_5_7, I8=>output_MAC_5_8, I9=>output_MAC_5_9, I10=>output_MAC_5_10, I11=>output_MAC_5_11, I12=>output_MAC_5_12, I13=>output_MAC_5_13, I14=>output_MAC_5_14, I15=>output_MAC_5_15, I16=>output_MAC_5_16, I17=>output_MAC_5_17, I18=>output_MAC_5_18, I19=>output_MAC_5_19, I20=>output_MAC_5_20, I21=>output_MAC_5_21, I22=>output_MAC_5_22, I23=>output_MAC_5_23, I24=>output_MAC_5_24, I25=>output_MAC_5_25, I26=>output_MAC_5_26, I27=>output_MAC_5_27, I28=>output_MAC_5_28, I29=>output_MAC_5_29, I30=>output_MAC_5_30, I31=>output_MAC_5_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_5);

	mux_row_6: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_6_0, I1=>output_MAC_6_1, I2=>output_MAC_6_2, I3=>output_MAC_6_3, I4=>output_MAC_6_4, I5=>output_MAC_6_5, I6=>output_MAC_6_6, I7=>output_MAC_6_7, I8=>output_MAC_6_8, I9=>output_MAC_6_9, I10=>output_MAC_6_10, I11=>output_MAC_6_11, I12=>output_MAC_6_12, I13=>output_MAC_6_13, I14=>output_MAC_6_14, I15=>output_MAC_6_15, I16=>output_MAC_6_16, I17=>output_MAC_6_17, I18=>output_MAC_6_18, I19=>output_MAC_6_19, I20=>output_MAC_6_20, I21=>output_MAC_6_21, I22=>output_MAC_6_22, I23=>output_MAC_6_23, I24=>output_MAC_6_24, I25=>output_MAC_6_25, I26=>output_MAC_6_26, I27=>output_MAC_6_27, I28=>output_MAC_6_28, I29=>output_MAC_6_29, I30=>output_MAC_6_30, I31=>output_MAC_6_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_6);

	mux_row_7: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_7_0, I1=>output_MAC_7_1, I2=>output_MAC_7_2, I3=>output_MAC_7_3, I4=>output_MAC_7_4, I5=>output_MAC_7_5, I6=>output_MAC_7_6, I7=>output_MAC_7_7, I8=>output_MAC_7_8, I9=>output_MAC_7_9, I10=>output_MAC_7_10, I11=>output_MAC_7_11, I12=>output_MAC_7_12, I13=>output_MAC_7_13, I14=>output_MAC_7_14, I15=>output_MAC_7_15, I16=>output_MAC_7_16, I17=>output_MAC_7_17, I18=>output_MAC_7_18, I19=>output_MAC_7_19, I20=>output_MAC_7_20, I21=>output_MAC_7_21, I22=>output_MAC_7_22, I23=>output_MAC_7_23, I24=>output_MAC_7_24, I25=>output_MAC_7_25, I26=>output_MAC_7_26, I27=>output_MAC_7_27, I28=>output_MAC_7_28, I29=>output_MAC_7_29, I30=>output_MAC_7_30, I31=>output_MAC_7_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_7);

	mux_row_8: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_8_0, I1=>output_MAC_8_1, I2=>output_MAC_8_2, I3=>output_MAC_8_3, I4=>output_MAC_8_4, I5=>output_MAC_8_5, I6=>output_MAC_8_6, I7=>output_MAC_8_7, I8=>output_MAC_8_8, I9=>output_MAC_8_9, I10=>output_MAC_8_10, I11=>output_MAC_8_11, I12=>output_MAC_8_12, I13=>output_MAC_8_13, I14=>output_MAC_8_14, I15=>output_MAC_8_15, I16=>output_MAC_8_16, I17=>output_MAC_8_17, I18=>output_MAC_8_18, I19=>output_MAC_8_19, I20=>output_MAC_8_20, I21=>output_MAC_8_21, I22=>output_MAC_8_22, I23=>output_MAC_8_23, I24=>output_MAC_8_24, I25=>output_MAC_8_25, I26=>output_MAC_8_26, I27=>output_MAC_8_27, I28=>output_MAC_8_28, I29=>output_MAC_8_29, I30=>output_MAC_8_30, I31=>output_MAC_8_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_8);

	mux_row_9: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_9_0, I1=>output_MAC_9_1, I2=>output_MAC_9_2, I3=>output_MAC_9_3, I4=>output_MAC_9_4, I5=>output_MAC_9_5, I6=>output_MAC_9_6, I7=>output_MAC_9_7, I8=>output_MAC_9_8, I9=>output_MAC_9_9, I10=>output_MAC_9_10, I11=>output_MAC_9_11, I12=>output_MAC_9_12, I13=>output_MAC_9_13, I14=>output_MAC_9_14, I15=>output_MAC_9_15, I16=>output_MAC_9_16, I17=>output_MAC_9_17, I18=>output_MAC_9_18, I19=>output_MAC_9_19, I20=>output_MAC_9_20, I21=>output_MAC_9_21, I22=>output_MAC_9_22, I23=>output_MAC_9_23, I24=>output_MAC_9_24, I25=>output_MAC_9_25, I26=>output_MAC_9_26, I27=>output_MAC_9_27, I28=>output_MAC_9_28, I29=>output_MAC_9_29, I30=>output_MAC_9_30, I31=>output_MAC_9_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_9);

	mux_row_10: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_10_0, I1=>output_MAC_10_1, I2=>output_MAC_10_2, I3=>output_MAC_10_3, I4=>output_MAC_10_4, I5=>output_MAC_10_5, I6=>output_MAC_10_6, I7=>output_MAC_10_7, I8=>output_MAC_10_8, I9=>output_MAC_10_9, I10=>output_MAC_10_10, I11=>output_MAC_10_11, I12=>output_MAC_10_12, I13=>output_MAC_10_13, I14=>output_MAC_10_14, I15=>output_MAC_10_15, I16=>output_MAC_10_16, I17=>output_MAC_10_17, I18=>output_MAC_10_18, I19=>output_MAC_10_19, I20=>output_MAC_10_20, I21=>output_MAC_10_21, I22=>output_MAC_10_22, I23=>output_MAC_10_23, I24=>output_MAC_10_24, I25=>output_MAC_10_25, I26=>output_MAC_10_26, I27=>output_MAC_10_27, I28=>output_MAC_10_28, I29=>output_MAC_10_29, I30=>output_MAC_10_30, I31=>output_MAC_10_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_10);

	mux_row_11: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_11_0, I1=>output_MAC_11_1, I2=>output_MAC_11_2, I3=>output_MAC_11_3, I4=>output_MAC_11_4, I5=>output_MAC_11_5, I6=>output_MAC_11_6, I7=>output_MAC_11_7, I8=>output_MAC_11_8, I9=>output_MAC_11_9, I10=>output_MAC_11_10, I11=>output_MAC_11_11, I12=>output_MAC_11_12, I13=>output_MAC_11_13, I14=>output_MAC_11_14, I15=>output_MAC_11_15, I16=>output_MAC_11_16, I17=>output_MAC_11_17, I18=>output_MAC_11_18, I19=>output_MAC_11_19, I20=>output_MAC_11_20, I21=>output_MAC_11_21, I22=>output_MAC_11_22, I23=>output_MAC_11_23, I24=>output_MAC_11_24, I25=>output_MAC_11_25, I26=>output_MAC_11_26, I27=>output_MAC_11_27, I28=>output_MAC_11_28, I29=>output_MAC_11_29, I30=>output_MAC_11_30, I31=>output_MAC_11_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_11);

	mux_row_12: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_12_0, I1=>output_MAC_12_1, I2=>output_MAC_12_2, I3=>output_MAC_12_3, I4=>output_MAC_12_4, I5=>output_MAC_12_5, I6=>output_MAC_12_6, I7=>output_MAC_12_7, I8=>output_MAC_12_8, I9=>output_MAC_12_9, I10=>output_MAC_12_10, I11=>output_MAC_12_11, I12=>output_MAC_12_12, I13=>output_MAC_12_13, I14=>output_MAC_12_14, I15=>output_MAC_12_15, I16=>output_MAC_12_16, I17=>output_MAC_12_17, I18=>output_MAC_12_18, I19=>output_MAC_12_19, I20=>output_MAC_12_20, I21=>output_MAC_12_21, I22=>output_MAC_12_22, I23=>output_MAC_12_23, I24=>output_MAC_12_24, I25=>output_MAC_12_25, I26=>output_MAC_12_26, I27=>output_MAC_12_27, I28=>output_MAC_12_28, I29=>output_MAC_12_29, I30=>output_MAC_12_30, I31=>output_MAC_12_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_12);

	mux_row_13: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_13_0, I1=>output_MAC_13_1, I2=>output_MAC_13_2, I3=>output_MAC_13_3, I4=>output_MAC_13_4, I5=>output_MAC_13_5, I6=>output_MAC_13_6, I7=>output_MAC_13_7, I8=>output_MAC_13_8, I9=>output_MAC_13_9, I10=>output_MAC_13_10, I11=>output_MAC_13_11, I12=>output_MAC_13_12, I13=>output_MAC_13_13, I14=>output_MAC_13_14, I15=>output_MAC_13_15, I16=>output_MAC_13_16, I17=>output_MAC_13_17, I18=>output_MAC_13_18, I19=>output_MAC_13_19, I20=>output_MAC_13_20, I21=>output_MAC_13_21, I22=>output_MAC_13_22, I23=>output_MAC_13_23, I24=>output_MAC_13_24, I25=>output_MAC_13_25, I26=>output_MAC_13_26, I27=>output_MAC_13_27, I28=>output_MAC_13_28, I29=>output_MAC_13_29, I30=>output_MAC_13_30, I31=>output_MAC_13_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_13);

	mux_row_14: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_14_0, I1=>output_MAC_14_1, I2=>output_MAC_14_2, I3=>output_MAC_14_3, I4=>output_MAC_14_4, I5=>output_MAC_14_5, I6=>output_MAC_14_6, I7=>output_MAC_14_7, I8=>output_MAC_14_8, I9=>output_MAC_14_9, I10=>output_MAC_14_10, I11=>output_MAC_14_11, I12=>output_MAC_14_12, I13=>output_MAC_14_13, I14=>output_MAC_14_14, I15=>output_MAC_14_15, I16=>output_MAC_14_16, I17=>output_MAC_14_17, I18=>output_MAC_14_18, I19=>output_MAC_14_19, I20=>output_MAC_14_20, I21=>output_MAC_14_21, I22=>output_MAC_14_22, I23=>output_MAC_14_23, I24=>output_MAC_14_24, I25=>output_MAC_14_25, I26=>output_MAC_14_26, I27=>output_MAC_14_27, I28=>output_MAC_14_28, I29=>output_MAC_14_29, I30=>output_MAC_14_30, I31=>output_MAC_14_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_14);

	mux_row_15: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_15_0, I1=>output_MAC_15_1, I2=>output_MAC_15_2, I3=>output_MAC_15_3, I4=>output_MAC_15_4, I5=>output_MAC_15_5, I6=>output_MAC_15_6, I7=>output_MAC_15_7, I8=>output_MAC_15_8, I9=>output_MAC_15_9, I10=>output_MAC_15_10, I11=>output_MAC_15_11, I12=>output_MAC_15_12, I13=>output_MAC_15_13, I14=>output_MAC_15_14, I15=>output_MAC_15_15, I16=>output_MAC_15_16, I17=>output_MAC_15_17, I18=>output_MAC_15_18, I19=>output_MAC_15_19, I20=>output_MAC_15_20, I21=>output_MAC_15_21, I22=>output_MAC_15_22, I23=>output_MAC_15_23, I24=>output_MAC_15_24, I25=>output_MAC_15_25, I26=>output_MAC_15_26, I27=>output_MAC_15_27, I28=>output_MAC_15_28, I29=>output_MAC_15_29, I30=>output_MAC_15_30, I31=>output_MAC_15_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_15);

	mux_row_16: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_16_0, I1=>output_MAC_16_1, I2=>output_MAC_16_2, I3=>output_MAC_16_3, I4=>output_MAC_16_4, I5=>output_MAC_16_5, I6=>output_MAC_16_6, I7=>output_MAC_16_7, I8=>output_MAC_16_8, I9=>output_MAC_16_9, I10=>output_MAC_16_10, I11=>output_MAC_16_11, I12=>output_MAC_16_12, I13=>output_MAC_16_13, I14=>output_MAC_16_14, I15=>output_MAC_16_15, I16=>output_MAC_16_16, I17=>output_MAC_16_17, I18=>output_MAC_16_18, I19=>output_MAC_16_19, I20=>output_MAC_16_20, I21=>output_MAC_16_21, I22=>output_MAC_16_22, I23=>output_MAC_16_23, I24=>output_MAC_16_24, I25=>output_MAC_16_25, I26=>output_MAC_16_26, I27=>output_MAC_16_27, I28=>output_MAC_16_28, I29=>output_MAC_16_29, I30=>output_MAC_16_30, I31=>output_MAC_16_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_16);

	mux_row_17: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_17_0, I1=>output_MAC_17_1, I2=>output_MAC_17_2, I3=>output_MAC_17_3, I4=>output_MAC_17_4, I5=>output_MAC_17_5, I6=>output_MAC_17_6, I7=>output_MAC_17_7, I8=>output_MAC_17_8, I9=>output_MAC_17_9, I10=>output_MAC_17_10, I11=>output_MAC_17_11, I12=>output_MAC_17_12, I13=>output_MAC_17_13, I14=>output_MAC_17_14, I15=>output_MAC_17_15, I16=>output_MAC_17_16, I17=>output_MAC_17_17, I18=>output_MAC_17_18, I19=>output_MAC_17_19, I20=>output_MAC_17_20, I21=>output_MAC_17_21, I22=>output_MAC_17_22, I23=>output_MAC_17_23, I24=>output_MAC_17_24, I25=>output_MAC_17_25, I26=>output_MAC_17_26, I27=>output_MAC_17_27, I28=>output_MAC_17_28, I29=>output_MAC_17_29, I30=>output_MAC_17_30, I31=>output_MAC_17_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_17);

	mux_row_18: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_18_0, I1=>output_MAC_18_1, I2=>output_MAC_18_2, I3=>output_MAC_18_3, I4=>output_MAC_18_4, I5=>output_MAC_18_5, I6=>output_MAC_18_6, I7=>output_MAC_18_7, I8=>output_MAC_18_8, I9=>output_MAC_18_9, I10=>output_MAC_18_10, I11=>output_MAC_18_11, I12=>output_MAC_18_12, I13=>output_MAC_18_13, I14=>output_MAC_18_14, I15=>output_MAC_18_15, I16=>output_MAC_18_16, I17=>output_MAC_18_17, I18=>output_MAC_18_18, I19=>output_MAC_18_19, I20=>output_MAC_18_20, I21=>output_MAC_18_21, I22=>output_MAC_18_22, I23=>output_MAC_18_23, I24=>output_MAC_18_24, I25=>output_MAC_18_25, I26=>output_MAC_18_26, I27=>output_MAC_18_27, I28=>output_MAC_18_28, I29=>output_MAC_18_29, I30=>output_MAC_18_30, I31=>output_MAC_18_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_18);

	mux_row_19: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_19_0, I1=>output_MAC_19_1, I2=>output_MAC_19_2, I3=>output_MAC_19_3, I4=>output_MAC_19_4, I5=>output_MAC_19_5, I6=>output_MAC_19_6, I7=>output_MAC_19_7, I8=>output_MAC_19_8, I9=>output_MAC_19_9, I10=>output_MAC_19_10, I11=>output_MAC_19_11, I12=>output_MAC_19_12, I13=>output_MAC_19_13, I14=>output_MAC_19_14, I15=>output_MAC_19_15, I16=>output_MAC_19_16, I17=>output_MAC_19_17, I18=>output_MAC_19_18, I19=>output_MAC_19_19, I20=>output_MAC_19_20, I21=>output_MAC_19_21, I22=>output_MAC_19_22, I23=>output_MAC_19_23, I24=>output_MAC_19_24, I25=>output_MAC_19_25, I26=>output_MAC_19_26, I27=>output_MAC_19_27, I28=>output_MAC_19_28, I29=>output_MAC_19_29, I30=>output_MAC_19_30, I31=>output_MAC_19_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_19);

	mux_row_20: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_20_0, I1=>output_MAC_20_1, I2=>output_MAC_20_2, I3=>output_MAC_20_3, I4=>output_MAC_20_4, I5=>output_MAC_20_5, I6=>output_MAC_20_6, I7=>output_MAC_20_7, I8=>output_MAC_20_8, I9=>output_MAC_20_9, I10=>output_MAC_20_10, I11=>output_MAC_20_11, I12=>output_MAC_20_12, I13=>output_MAC_20_13, I14=>output_MAC_20_14, I15=>output_MAC_20_15, I16=>output_MAC_20_16, I17=>output_MAC_20_17, I18=>output_MAC_20_18, I19=>output_MAC_20_19, I20=>output_MAC_20_20, I21=>output_MAC_20_21, I22=>output_MAC_20_22, I23=>output_MAC_20_23, I24=>output_MAC_20_24, I25=>output_MAC_20_25, I26=>output_MAC_20_26, I27=>output_MAC_20_27, I28=>output_MAC_20_28, I29=>output_MAC_20_29, I30=>output_MAC_20_30, I31=>output_MAC_20_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_20);

	mux_row_21: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_21_0, I1=>output_MAC_21_1, I2=>output_MAC_21_2, I3=>output_MAC_21_3, I4=>output_MAC_21_4, I5=>output_MAC_21_5, I6=>output_MAC_21_6, I7=>output_MAC_21_7, I8=>output_MAC_21_8, I9=>output_MAC_21_9, I10=>output_MAC_21_10, I11=>output_MAC_21_11, I12=>output_MAC_21_12, I13=>output_MAC_21_13, I14=>output_MAC_21_14, I15=>output_MAC_21_15, I16=>output_MAC_21_16, I17=>output_MAC_21_17, I18=>output_MAC_21_18, I19=>output_MAC_21_19, I20=>output_MAC_21_20, I21=>output_MAC_21_21, I22=>output_MAC_21_22, I23=>output_MAC_21_23, I24=>output_MAC_21_24, I25=>output_MAC_21_25, I26=>output_MAC_21_26, I27=>output_MAC_21_27, I28=>output_MAC_21_28, I29=>output_MAC_21_29, I30=>output_MAC_21_30, I31=>output_MAC_21_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_21);

	mux_row_22: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_22_0, I1=>output_MAC_22_1, I2=>output_MAC_22_2, I3=>output_MAC_22_3, I4=>output_MAC_22_4, I5=>output_MAC_22_5, I6=>output_MAC_22_6, I7=>output_MAC_22_7, I8=>output_MAC_22_8, I9=>output_MAC_22_9, I10=>output_MAC_22_10, I11=>output_MAC_22_11, I12=>output_MAC_22_12, I13=>output_MAC_22_13, I14=>output_MAC_22_14, I15=>output_MAC_22_15, I16=>output_MAC_22_16, I17=>output_MAC_22_17, I18=>output_MAC_22_18, I19=>output_MAC_22_19, I20=>output_MAC_22_20, I21=>output_MAC_22_21, I22=>output_MAC_22_22, I23=>output_MAC_22_23, I24=>output_MAC_22_24, I25=>output_MAC_22_25, I26=>output_MAC_22_26, I27=>output_MAC_22_27, I28=>output_MAC_22_28, I29=>output_MAC_22_29, I30=>output_MAC_22_30, I31=>output_MAC_22_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_22);

	mux_row_23: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_23_0, I1=>output_MAC_23_1, I2=>output_MAC_23_2, I3=>output_MAC_23_3, I4=>output_MAC_23_4, I5=>output_MAC_23_5, I6=>output_MAC_23_6, I7=>output_MAC_23_7, I8=>output_MAC_23_8, I9=>output_MAC_23_9, I10=>output_MAC_23_10, I11=>output_MAC_23_11, I12=>output_MAC_23_12, I13=>output_MAC_23_13, I14=>output_MAC_23_14, I15=>output_MAC_23_15, I16=>output_MAC_23_16, I17=>output_MAC_23_17, I18=>output_MAC_23_18, I19=>output_MAC_23_19, I20=>output_MAC_23_20, I21=>output_MAC_23_21, I22=>output_MAC_23_22, I23=>output_MAC_23_23, I24=>output_MAC_23_24, I25=>output_MAC_23_25, I26=>output_MAC_23_26, I27=>output_MAC_23_27, I28=>output_MAC_23_28, I29=>output_MAC_23_29, I30=>output_MAC_23_30, I31=>output_MAC_23_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_23);

	mux_row_24: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_24_0, I1=>output_MAC_24_1, I2=>output_MAC_24_2, I3=>output_MAC_24_3, I4=>output_MAC_24_4, I5=>output_MAC_24_5, I6=>output_MAC_24_6, I7=>output_MAC_24_7, I8=>output_MAC_24_8, I9=>output_MAC_24_9, I10=>output_MAC_24_10, I11=>output_MAC_24_11, I12=>output_MAC_24_12, I13=>output_MAC_24_13, I14=>output_MAC_24_14, I15=>output_MAC_24_15, I16=>output_MAC_24_16, I17=>output_MAC_24_17, I18=>output_MAC_24_18, I19=>output_MAC_24_19, I20=>output_MAC_24_20, I21=>output_MAC_24_21, I22=>output_MAC_24_22, I23=>output_MAC_24_23, I24=>output_MAC_24_24, I25=>output_MAC_24_25, I26=>output_MAC_24_26, I27=>output_MAC_24_27, I28=>output_MAC_24_28, I29=>output_MAC_24_29, I30=>output_MAC_24_30, I31=>output_MAC_24_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_24);

	mux_row_25: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_25_0, I1=>output_MAC_25_1, I2=>output_MAC_25_2, I3=>output_MAC_25_3, I4=>output_MAC_25_4, I5=>output_MAC_25_5, I6=>output_MAC_25_6, I7=>output_MAC_25_7, I8=>output_MAC_25_8, I9=>output_MAC_25_9, I10=>output_MAC_25_10, I11=>output_MAC_25_11, I12=>output_MAC_25_12, I13=>output_MAC_25_13, I14=>output_MAC_25_14, I15=>output_MAC_25_15, I16=>output_MAC_25_16, I17=>output_MAC_25_17, I18=>output_MAC_25_18, I19=>output_MAC_25_19, I20=>output_MAC_25_20, I21=>output_MAC_25_21, I22=>output_MAC_25_22, I23=>output_MAC_25_23, I24=>output_MAC_25_24, I25=>output_MAC_25_25, I26=>output_MAC_25_26, I27=>output_MAC_25_27, I28=>output_MAC_25_28, I29=>output_MAC_25_29, I30=>output_MAC_25_30, I31=>output_MAC_25_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_25);

	mux_row_26: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_26_0, I1=>output_MAC_26_1, I2=>output_MAC_26_2, I3=>output_MAC_26_3, I4=>output_MAC_26_4, I5=>output_MAC_26_5, I6=>output_MAC_26_6, I7=>output_MAC_26_7, I8=>output_MAC_26_8, I9=>output_MAC_26_9, I10=>output_MAC_26_10, I11=>output_MAC_26_11, I12=>output_MAC_26_12, I13=>output_MAC_26_13, I14=>output_MAC_26_14, I15=>output_MAC_26_15, I16=>output_MAC_26_16, I17=>output_MAC_26_17, I18=>output_MAC_26_18, I19=>output_MAC_26_19, I20=>output_MAC_26_20, I21=>output_MAC_26_21, I22=>output_MAC_26_22, I23=>output_MAC_26_23, I24=>output_MAC_26_24, I25=>output_MAC_26_25, I26=>output_MAC_26_26, I27=>output_MAC_26_27, I28=>output_MAC_26_28, I29=>output_MAC_26_29, I30=>output_MAC_26_30, I31=>output_MAC_26_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_26);

	mux_row_27: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_27_0, I1=>output_MAC_27_1, I2=>output_MAC_27_2, I3=>output_MAC_27_3, I4=>output_MAC_27_4, I5=>output_MAC_27_5, I6=>output_MAC_27_6, I7=>output_MAC_27_7, I8=>output_MAC_27_8, I9=>output_MAC_27_9, I10=>output_MAC_27_10, I11=>output_MAC_27_11, I12=>output_MAC_27_12, I13=>output_MAC_27_13, I14=>output_MAC_27_14, I15=>output_MAC_27_15, I16=>output_MAC_27_16, I17=>output_MAC_27_17, I18=>output_MAC_27_18, I19=>output_MAC_27_19, I20=>output_MAC_27_20, I21=>output_MAC_27_21, I22=>output_MAC_27_22, I23=>output_MAC_27_23, I24=>output_MAC_27_24, I25=>output_MAC_27_25, I26=>output_MAC_27_26, I27=>output_MAC_27_27, I28=>output_MAC_27_28, I29=>output_MAC_27_29, I30=>output_MAC_27_30, I31=>output_MAC_27_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_27);

	mux_row_28: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_28_0, I1=>output_MAC_28_1, I2=>output_MAC_28_2, I3=>output_MAC_28_3, I4=>output_MAC_28_4, I5=>output_MAC_28_5, I6=>output_MAC_28_6, I7=>output_MAC_28_7, I8=>output_MAC_28_8, I9=>output_MAC_28_9, I10=>output_MAC_28_10, I11=>output_MAC_28_11, I12=>output_MAC_28_12, I13=>output_MAC_28_13, I14=>output_MAC_28_14, I15=>output_MAC_28_15, I16=>output_MAC_28_16, I17=>output_MAC_28_17, I18=>output_MAC_28_18, I19=>output_MAC_28_19, I20=>output_MAC_28_20, I21=>output_MAC_28_21, I22=>output_MAC_28_22, I23=>output_MAC_28_23, I24=>output_MAC_28_24, I25=>output_MAC_28_25, I26=>output_MAC_28_26, I27=>output_MAC_28_27, I28=>output_MAC_28_28, I29=>output_MAC_28_29, I30=>output_MAC_28_30, I31=>output_MAC_28_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_28);

	mux_row_29: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_29_0, I1=>output_MAC_29_1, I2=>output_MAC_29_2, I3=>output_MAC_29_3, I4=>output_MAC_29_4, I5=>output_MAC_29_5, I6=>output_MAC_29_6, I7=>output_MAC_29_7, I8=>output_MAC_29_8, I9=>output_MAC_29_9, I10=>output_MAC_29_10, I11=>output_MAC_29_11, I12=>output_MAC_29_12, I13=>output_MAC_29_13, I14=>output_MAC_29_14, I15=>output_MAC_29_15, I16=>output_MAC_29_16, I17=>output_MAC_29_17, I18=>output_MAC_29_18, I19=>output_MAC_29_19, I20=>output_MAC_29_20, I21=>output_MAC_29_21, I22=>output_MAC_29_22, I23=>output_MAC_29_23, I24=>output_MAC_29_24, I25=>output_MAC_29_25, I26=>output_MAC_29_26, I27=>output_MAC_29_27, I28=>output_MAC_29_28, I29=>output_MAC_29_29, I30=>output_MAC_29_30, I31=>output_MAC_29_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_29);

	mux_row_30: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_30_0, I1=>output_MAC_30_1, I2=>output_MAC_30_2, I3=>output_MAC_30_3, I4=>output_MAC_30_4, I5=>output_MAC_30_5, I6=>output_MAC_30_6, I7=>output_MAC_30_7, I8=>output_MAC_30_8, I9=>output_MAC_30_9, I10=>output_MAC_30_10, I11=>output_MAC_30_11, I12=>output_MAC_30_12, I13=>output_MAC_30_13, I14=>output_MAC_30_14, I15=>output_MAC_30_15, I16=>output_MAC_30_16, I17=>output_MAC_30_17, I18=>output_MAC_30_18, I19=>output_MAC_30_19, I20=>output_MAC_30_20, I21=>output_MAC_30_21, I22=>output_MAC_30_22, I23=>output_MAC_30_23, I24=>output_MAC_30_24, I25=>output_MAC_30_25, I26=>output_MAC_30_26, I27=>output_MAC_30_27, I28=>output_MAC_30_28, I29=>output_MAC_30_29, I30=>output_MAC_30_30, I31=>output_MAC_30_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_30);

	mux_row_31: mux_32to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_31_0, I1=>output_MAC_31_1, I2=>output_MAC_31_2, I3=>output_MAC_31_3, I4=>output_MAC_31_4, I5=>output_MAC_31_5, I6=>output_MAC_31_6, I7=>output_MAC_31_7, I8=>output_MAC_31_8, I9=>output_MAC_31_9, I10=>output_MAC_31_10, I11=>output_MAC_31_11, I12=>output_MAC_31_12, I13=>output_MAC_31_13, I14=>output_MAC_31_14, I15=>output_MAC_31_15, I16=>output_MAC_31_16, I17=>output_MAC_31_17, I18=>output_MAC_31_18, I19=>output_MAC_31_19, I20=>output_MAC_31_20, I21=>output_MAC_31_21, I22=>output_MAC_31_22, I23=>output_MAC_31_23, I24=>output_MAC_31_24, I25=>output_MAC_31_25, I26=>output_MAC_31_26, I27=>output_MAC_31_27, I28=>output_MAC_31_28, I29=>output_MAC_31_29, I30=>output_MAC_31_30, I31=>output_MAC_31_31, 
		SEL_mux=>reg_SEL_mux, O=>reg_output_row_31);

	output_row_0_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_0, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_0);
	output_row_1_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_1, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_1);
	output_row_2_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_2, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_2);
	output_row_3_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_3, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_3);
	output_row_4_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_4, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_4);
	output_row_5_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_5, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_5);
	output_row_6_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_6, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_6);
	output_row_7_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_7, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_7);
	output_row_8_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_8, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_8);
	output_row_9_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_9, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_9);
	output_row_10_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_10, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_10);
	output_row_11_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_11, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_11);
	output_row_12_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_12, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_12);
	output_row_13_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_13, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_13);
	output_row_14_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_14, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_14);
	output_row_15_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_15, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_15);
	output_row_16_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_16, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_16);
	output_row_17_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_17, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_17);
	output_row_18_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_18, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_18);
	output_row_19_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_19, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_19);
	output_row_20_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_20, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_20);
	output_row_21_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_21, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_21);
	output_row_22_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_22, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_22);
	output_row_23_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_23, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_23);
	output_row_24_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_24, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_24);
	output_row_25_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_25, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_25);
	output_row_26_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_26, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_26);
	output_row_27_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_27, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_27);
	output_row_28_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_28, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_28);
	output_row_29_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_29, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_29);
	output_row_30_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_30, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_30);
	output_row_31_reg: regnbit GENERIC MAP(N=>32)
		PORT MAP(D=>reg_output_row_31, CLK=>CLK, RST_n=>RST_n, ENABLE=>'1', Q=>output_row_31);

END behaviour;
