
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MAC_8x768_8 IS
PORT (input_row_0, input_row_1, input_row_2, input_row_3, input_row_4, input_row_5, input_row_6, input_row_7: IN STD_LOGIC_VECTOR(7 downto 0);
	input_col_0, input_col_1, input_col_2, input_col_3, input_col_4, input_col_5, input_col_6, input_col_7, input_col_8, input_col_9, 
	input_col_10, input_col_11, input_col_12, input_col_13, input_col_14, input_col_15, input_col_16, input_col_17, input_col_18, input_col_19, 
	input_col_20, input_col_21, input_col_22, input_col_23, input_col_24, input_col_25, input_col_26, input_col_27, input_col_28, input_col_29, 
	input_col_30, input_col_31, input_col_32, input_col_33, input_col_34, input_col_35, input_col_36, input_col_37, input_col_38, input_col_39, 
	input_col_40, input_col_41, input_col_42, input_col_43, input_col_44, input_col_45, input_col_46, input_col_47, input_col_48, input_col_49, 
	input_col_50, input_col_51, input_col_52, input_col_53, input_col_54, input_col_55, input_col_56, input_col_57, input_col_58, input_col_59, 
	input_col_60, input_col_61, input_col_62, input_col_63, input_col_64, input_col_65, input_col_66, input_col_67, input_col_68, input_col_69, 
	input_col_70, input_col_71, input_col_72, input_col_73, input_col_74, input_col_75, input_col_76, input_col_77, input_col_78, input_col_79, 
	input_col_80, input_col_81, input_col_82, input_col_83, input_col_84, input_col_85, input_col_86, input_col_87, input_col_88, input_col_89, 
	input_col_90, input_col_91, input_col_92, input_col_93, input_col_94, input_col_95, input_col_96, input_col_97, input_col_98, input_col_99, 
	input_col_100, input_col_101, input_col_102, input_col_103, input_col_104, input_col_105, input_col_106, input_col_107, input_col_108, input_col_109, 
	input_col_110, input_col_111, input_col_112, input_col_113, input_col_114, input_col_115, input_col_116, input_col_117, input_col_118, input_col_119, 
	input_col_120, input_col_121, input_col_122, input_col_123, input_col_124, input_col_125, input_col_126, input_col_127, input_col_128, input_col_129, 
	input_col_130, input_col_131, input_col_132, input_col_133, input_col_134, input_col_135, input_col_136, input_col_137, input_col_138, input_col_139, 
	input_col_140, input_col_141, input_col_142, input_col_143, input_col_144, input_col_145, input_col_146, input_col_147, input_col_148, input_col_149, 
	input_col_150, input_col_151, input_col_152, input_col_153, input_col_154, input_col_155, input_col_156, input_col_157, input_col_158, input_col_159, 
	input_col_160, input_col_161, input_col_162, input_col_163, input_col_164, input_col_165, input_col_166, input_col_167, input_col_168, input_col_169, 
	input_col_170, input_col_171, input_col_172, input_col_173, input_col_174, input_col_175, input_col_176, input_col_177, input_col_178, input_col_179, 
	input_col_180, input_col_181, input_col_182, input_col_183, input_col_184, input_col_185, input_col_186, input_col_187, input_col_188, input_col_189, 
	input_col_190, input_col_191, input_col_192, input_col_193, input_col_194, input_col_195, input_col_196, input_col_197, input_col_198, input_col_199, 
	input_col_200, input_col_201, input_col_202, input_col_203, input_col_204, input_col_205, input_col_206, input_col_207, input_col_208, input_col_209, 
	input_col_210, input_col_211, input_col_212, input_col_213, input_col_214, input_col_215, input_col_216, input_col_217, input_col_218, input_col_219, 
	input_col_220, input_col_221, input_col_222, input_col_223, input_col_224, input_col_225, input_col_226, input_col_227, input_col_228, input_col_229, 
	input_col_230, input_col_231, input_col_232, input_col_233, input_col_234, input_col_235, input_col_236, input_col_237, input_col_238, input_col_239, 
	input_col_240, input_col_241, input_col_242, input_col_243, input_col_244, input_col_245, input_col_246, input_col_247, input_col_248, input_col_249, 
	input_col_250, input_col_251, input_col_252, input_col_253, input_col_254, input_col_255, input_col_256, input_col_257, input_col_258, input_col_259, 
	input_col_260, input_col_261, input_col_262, input_col_263, input_col_264, input_col_265, input_col_266, input_col_267, input_col_268, input_col_269, 
	input_col_270, input_col_271, input_col_272, input_col_273, input_col_274, input_col_275, input_col_276, input_col_277, input_col_278, input_col_279, 
	input_col_280, input_col_281, input_col_282, input_col_283, input_col_284, input_col_285, input_col_286, input_col_287, input_col_288, input_col_289, 
	input_col_290, input_col_291, input_col_292, input_col_293, input_col_294, input_col_295, input_col_296, input_col_297, input_col_298, input_col_299, 
	input_col_300, input_col_301, input_col_302, input_col_303, input_col_304, input_col_305, input_col_306, input_col_307, input_col_308, input_col_309, 
	input_col_310, input_col_311, input_col_312, input_col_313, input_col_314, input_col_315, input_col_316, input_col_317, input_col_318, input_col_319, 
	input_col_320, input_col_321, input_col_322, input_col_323, input_col_324, input_col_325, input_col_326, input_col_327, input_col_328, input_col_329, 
	input_col_330, input_col_331, input_col_332, input_col_333, input_col_334, input_col_335, input_col_336, input_col_337, input_col_338, input_col_339, 
	input_col_340, input_col_341, input_col_342, input_col_343, input_col_344, input_col_345, input_col_346, input_col_347, input_col_348, input_col_349, 
	input_col_350, input_col_351, input_col_352, input_col_353, input_col_354, input_col_355, input_col_356, input_col_357, input_col_358, input_col_359, 
	input_col_360, input_col_361, input_col_362, input_col_363, input_col_364, input_col_365, input_col_366, input_col_367, input_col_368, input_col_369, 
	input_col_370, input_col_371, input_col_372, input_col_373, input_col_374, input_col_375, input_col_376, input_col_377, input_col_378, input_col_379, 
	input_col_380, input_col_381, input_col_382, input_col_383, input_col_384, input_col_385, input_col_386, input_col_387, input_col_388, input_col_389, 
	input_col_390, input_col_391, input_col_392, input_col_393, input_col_394, input_col_395, input_col_396, input_col_397, input_col_398, input_col_399, 
	input_col_400, input_col_401, input_col_402, input_col_403, input_col_404, input_col_405, input_col_406, input_col_407, input_col_408, input_col_409, 
	input_col_410, input_col_411, input_col_412, input_col_413, input_col_414, input_col_415, input_col_416, input_col_417, input_col_418, input_col_419, 
	input_col_420, input_col_421, input_col_422, input_col_423, input_col_424, input_col_425, input_col_426, input_col_427, input_col_428, input_col_429, 
	input_col_430, input_col_431, input_col_432, input_col_433, input_col_434, input_col_435, input_col_436, input_col_437, input_col_438, input_col_439, 
	input_col_440, input_col_441, input_col_442, input_col_443, input_col_444, input_col_445, input_col_446, input_col_447, input_col_448, input_col_449, 
	input_col_450, input_col_451, input_col_452, input_col_453, input_col_454, input_col_455, input_col_456, input_col_457, input_col_458, input_col_459, 
	input_col_460, input_col_461, input_col_462, input_col_463, input_col_464, input_col_465, input_col_466, input_col_467, input_col_468, input_col_469, 
	input_col_470, input_col_471, input_col_472, input_col_473, input_col_474, input_col_475, input_col_476, input_col_477, input_col_478, input_col_479, 
	input_col_480, input_col_481, input_col_482, input_col_483, input_col_484, input_col_485, input_col_486, input_col_487, input_col_488, input_col_489, 
	input_col_490, input_col_491, input_col_492, input_col_493, input_col_494, input_col_495, input_col_496, input_col_497, input_col_498, input_col_499, 
	input_col_500, input_col_501, input_col_502, input_col_503, input_col_504, input_col_505, input_col_506, input_col_507, input_col_508, input_col_509, 
	input_col_510, input_col_511, input_col_512, input_col_513, input_col_514, input_col_515, input_col_516, input_col_517, input_col_518, input_col_519, 
	input_col_520, input_col_521, input_col_522, input_col_523, input_col_524, input_col_525, input_col_526, input_col_527, input_col_528, input_col_529, 
	input_col_530, input_col_531, input_col_532, input_col_533, input_col_534, input_col_535, input_col_536, input_col_537, input_col_538, input_col_539, 
	input_col_540, input_col_541, input_col_542, input_col_543, input_col_544, input_col_545, input_col_546, input_col_547, input_col_548, input_col_549, 
	input_col_550, input_col_551, input_col_552, input_col_553, input_col_554, input_col_555, input_col_556, input_col_557, input_col_558, input_col_559, 
	input_col_560, input_col_561, input_col_562, input_col_563, input_col_564, input_col_565, input_col_566, input_col_567, input_col_568, input_col_569, 
	input_col_570, input_col_571, input_col_572, input_col_573, input_col_574, input_col_575, input_col_576, input_col_577, input_col_578, input_col_579, 
	input_col_580, input_col_581, input_col_582, input_col_583, input_col_584, input_col_585, input_col_586, input_col_587, input_col_588, input_col_589, 
	input_col_590, input_col_591, input_col_592, input_col_593, input_col_594, input_col_595, input_col_596, input_col_597, input_col_598, input_col_599, 
	input_col_600, input_col_601, input_col_602, input_col_603, input_col_604, input_col_605, input_col_606, input_col_607, input_col_608, input_col_609, 
	input_col_610, input_col_611, input_col_612, input_col_613, input_col_614, input_col_615, input_col_616, input_col_617, input_col_618, input_col_619, 
	input_col_620, input_col_621, input_col_622, input_col_623, input_col_624, input_col_625, input_col_626, input_col_627, input_col_628, input_col_629, 
	input_col_630, input_col_631, input_col_632, input_col_633, input_col_634, input_col_635, input_col_636, input_col_637, input_col_638, input_col_639, 
	input_col_640, input_col_641, input_col_642, input_col_643, input_col_644, input_col_645, input_col_646, input_col_647, input_col_648, input_col_649, 
	input_col_650, input_col_651, input_col_652, input_col_653, input_col_654, input_col_655, input_col_656, input_col_657, input_col_658, input_col_659, 
	input_col_660, input_col_661, input_col_662, input_col_663, input_col_664, input_col_665, input_col_666, input_col_667, input_col_668, input_col_669, 
	input_col_670, input_col_671, input_col_672, input_col_673, input_col_674, input_col_675, input_col_676, input_col_677, input_col_678, input_col_679, 
	input_col_680, input_col_681, input_col_682, input_col_683, input_col_684, input_col_685, input_col_686, input_col_687, input_col_688, input_col_689, 
	input_col_690, input_col_691, input_col_692, input_col_693, input_col_694, input_col_695, input_col_696, input_col_697, input_col_698, input_col_699, 
	input_col_700, input_col_701, input_col_702, input_col_703, input_col_704, input_col_705, input_col_706, input_col_707, input_col_708, input_col_709, 
	input_col_710, input_col_711, input_col_712, input_col_713, input_col_714, input_col_715, input_col_716, input_col_717, input_col_718, input_col_719, 
	input_col_720, input_col_721, input_col_722, input_col_723, input_col_724, input_col_725, input_col_726, input_col_727, input_col_728, input_col_729, 
	input_col_730, input_col_731, input_col_732, input_col_733, input_col_734, input_col_735, input_col_736, input_col_737, input_col_738, input_col_739, 
	input_col_740, input_col_741, input_col_742, input_col_743, input_col_744, input_col_745, input_col_746, input_col_747, input_col_748, input_col_749, 
	input_col_750, input_col_751, input_col_752, input_col_753, input_col_754, input_col_755, input_col_756, input_col_757, input_col_758, input_col_759, 
	input_col_760, input_col_761, input_col_762, input_col_763, input_col_764, input_col_765, input_col_766, input_col_767: IN STD_LOGIC_VECTOR(7 downto 0);
	SEL_mux: IN STD_LOGIC_VECTOR(9 downto 0);
	CLK, RST_n, ENABLE : IN STD_LOGIC;
	output_row_0, output_row_1, output_row_2, output_row_3, output_row_4, output_row_5, output_row_6, output_row_7: OUT STD_LOGIC_VECTOR(31 downto 0)
);
END MAC_8x768_8;

ARCHITECTURE behaviour OF  MAC_8x768_8 IS

	COMPONENT MAC IS
	GENERIC (data_size : POSITIVE := 2;
	 acc_size : POSITIVE := 16 );
	PORT( data_in_A, data_in_B  : IN STD_LOGIC_VECTOR(data_size-1 downto 0);
		CLK, RST_n, ENABLE 	: IN STD_LOGIC;
		data_out    			: OUT STD_LOGIC_VECTOR(acc_size-1 downto 0));
	END COMPONENT;

	COMPONENT mux_768to1_nbit IS
	GENERIC ( N : POSITIVE :=2);
	PORT(
		I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, 
		I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, 
		I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, 
		I30, I31, I32, I33, I34, I35, I36, I37, I38, I39, 
		I40, I41, I42, I43, I44, I45, I46, I47, I48, I49, 
		I50, I51, I52, I53, I54, I55, I56, I57, I58, I59, 
		I60, I61, I62, I63, I64, I65, I66, I67, I68, I69, 
		I70, I71, I72, I73, I74, I75, I76, I77, I78, I79, 
		I80, I81, I82, I83, I84, I85, I86, I87, I88, I89, 
		I90, I91, I92, I93, I94, I95, I96, I97, I98, I99, 
		I100, I101, I102, I103, I104, I105, I106, I107, I108, I109, 
		I110, I111, I112, I113, I114, I115, I116, I117, I118, I119, 
		I120, I121, I122, I123, I124, I125, I126, I127, I128, I129, 
		I130, I131, I132, I133, I134, I135, I136, I137, I138, I139, 
		I140, I141, I142, I143, I144, I145, I146, I147, I148, I149, 
		I150, I151, I152, I153, I154, I155, I156, I157, I158, I159, 
		I160, I161, I162, I163, I164, I165, I166, I167, I168, I169, 
		I170, I171, I172, I173, I174, I175, I176, I177, I178, I179, 
		I180, I181, I182, I183, I184, I185, I186, I187, I188, I189, 
		I190, I191, I192, I193, I194, I195, I196, I197, I198, I199, 
		I200, I201, I202, I203, I204, I205, I206, I207, I208, I209, 
		I210, I211, I212, I213, I214, I215, I216, I217, I218, I219, 
		I220, I221, I222, I223, I224, I225, I226, I227, I228, I229, 
		I230, I231, I232, I233, I234, I235, I236, I237, I238, I239, 
		I240, I241, I242, I243, I244, I245, I246, I247, I248, I249, 
		I250, I251, I252, I253, I254, I255, I256, I257, I258, I259, 
		I260, I261, I262, I263, I264, I265, I266, I267, I268, I269, 
		I270, I271, I272, I273, I274, I275, I276, I277, I278, I279, 
		I280, I281, I282, I283, I284, I285, I286, I287, I288, I289, 
		I290, I291, I292, I293, I294, I295, I296, I297, I298, I299, 
		I300, I301, I302, I303, I304, I305, I306, I307, I308, I309, 
		I310, I311, I312, I313, I314, I315, I316, I317, I318, I319, 
		I320, I321, I322, I323, I324, I325, I326, I327, I328, I329, 
		I330, I331, I332, I333, I334, I335, I336, I337, I338, I339, 
		I340, I341, I342, I343, I344, I345, I346, I347, I348, I349, 
		I350, I351, I352, I353, I354, I355, I356, I357, I358, I359, 
		I360, I361, I362, I363, I364, I365, I366, I367, I368, I369, 
		I370, I371, I372, I373, I374, I375, I376, I377, I378, I379, 
		I380, I381, I382, I383, I384, I385, I386, I387, I388, I389, 
		I390, I391, I392, I393, I394, I395, I396, I397, I398, I399, 
		I400, I401, I402, I403, I404, I405, I406, I407, I408, I409, 
		I410, I411, I412, I413, I414, I415, I416, I417, I418, I419, 
		I420, I421, I422, I423, I424, I425, I426, I427, I428, I429, 
		I430, I431, I432, I433, I434, I435, I436, I437, I438, I439, 
		I440, I441, I442, I443, I444, I445, I446, I447, I448, I449, 
		I450, I451, I452, I453, I454, I455, I456, I457, I458, I459, 
		I460, I461, I462, I463, I464, I465, I466, I467, I468, I469, 
		I470, I471, I472, I473, I474, I475, I476, I477, I478, I479, 
		I480, I481, I482, I483, I484, I485, I486, I487, I488, I489, 
		I490, I491, I492, I493, I494, I495, I496, I497, I498, I499, 
		I500, I501, I502, I503, I504, I505, I506, I507, I508, I509, 
		I510, I511, I512, I513, I514, I515, I516, I517, I518, I519, 
		I520, I521, I522, I523, I524, I525, I526, I527, I528, I529, 
		I530, I531, I532, I533, I534, I535, I536, I537, I538, I539, 
		I540, I541, I542, I543, I544, I545, I546, I547, I548, I549, 
		I550, I551, I552, I553, I554, I555, I556, I557, I558, I559, 
		I560, I561, I562, I563, I564, I565, I566, I567, I568, I569, 
		I570, I571, I572, I573, I574, I575, I576, I577, I578, I579, 
		I580, I581, I582, I583, I584, I585, I586, I587, I588, I589, 
		I590, I591, I592, I593, I594, I595, I596, I597, I598, I599, 
		I600, I601, I602, I603, I604, I605, I606, I607, I608, I609, 
		I610, I611, I612, I613, I614, I615, I616, I617, I618, I619, 
		I620, I621, I622, I623, I624, I625, I626, I627, I628, I629, 
		I630, I631, I632, I633, I634, I635, I636, I637, I638, I639, 
		I640, I641, I642, I643, I644, I645, I646, I647, I648, I649, 
		I650, I651, I652, I653, I654, I655, I656, I657, I658, I659, 
		I660, I661, I662, I663, I664, I665, I666, I667, I668, I669, 
		I670, I671, I672, I673, I674, I675, I676, I677, I678, I679, 
		I680, I681, I682, I683, I684, I685, I686, I687, I688, I689, 
		I690, I691, I692, I693, I694, I695, I696, I697, I698, I699, 
		I700, I701, I702, I703, I704, I705, I706, I707, I708, I709, 
		I710, I711, I712, I713, I714, I715, I716, I717, I718, I719, 
		I720, I721, I722, I723, I724, I725, I726, I727, I728, I729, 
		I730, I731, I732, I733, I734, I735, I736, I737, I738, I739, 
		I740, I741, I742, I743, I744, I745, I746, I747, I748, I749, 
		I750, I751, I752, I753, I754, I755, I756, I757, I758, I759, 
		I760, I761, I762, I763, I764, I765, I766, I767: IN STD_LOGIC_VECTOR(N-1 downto 0);
		SEL_mux  : IN STD_LOGIC_VECTOR(9 downto 0);
		O    : OUT STD_LOGIC_VECTOR(N-1 downto 0)
	);
	END COMPONENT;


	SIGNAL output_MAC_0_0, output_MAC_0_1, output_MAC_0_2, output_MAC_0_3, output_MAC_0_4, output_MAC_0_5, output_MAC_0_6, output_MAC_0_7, output_MAC_0_8, output_MAC_0_9, 
		output_MAC_0_10, output_MAC_0_11, output_MAC_0_12, output_MAC_0_13, output_MAC_0_14, output_MAC_0_15, output_MAC_0_16, output_MAC_0_17, output_MAC_0_18, output_MAC_0_19, 
		output_MAC_0_20, output_MAC_0_21, output_MAC_0_22, output_MAC_0_23, output_MAC_0_24, output_MAC_0_25, output_MAC_0_26, output_MAC_0_27, output_MAC_0_28, output_MAC_0_29, 
		output_MAC_0_30, output_MAC_0_31, output_MAC_0_32, output_MAC_0_33, output_MAC_0_34, output_MAC_0_35, output_MAC_0_36, output_MAC_0_37, output_MAC_0_38, output_MAC_0_39, 
		output_MAC_0_40, output_MAC_0_41, output_MAC_0_42, output_MAC_0_43, output_MAC_0_44, output_MAC_0_45, output_MAC_0_46, output_MAC_0_47, output_MAC_0_48, output_MAC_0_49, 
		output_MAC_0_50, output_MAC_0_51, output_MAC_0_52, output_MAC_0_53, output_MAC_0_54, output_MAC_0_55, output_MAC_0_56, output_MAC_0_57, output_MAC_0_58, output_MAC_0_59, 
		output_MAC_0_60, output_MAC_0_61, output_MAC_0_62, output_MAC_0_63, output_MAC_0_64, output_MAC_0_65, output_MAC_0_66, output_MAC_0_67, output_MAC_0_68, output_MAC_0_69, 
		output_MAC_0_70, output_MAC_0_71, output_MAC_0_72, output_MAC_0_73, output_MAC_0_74, output_MAC_0_75, output_MAC_0_76, output_MAC_0_77, output_MAC_0_78, output_MAC_0_79, 
		output_MAC_0_80, output_MAC_0_81, output_MAC_0_82, output_MAC_0_83, output_MAC_0_84, output_MAC_0_85, output_MAC_0_86, output_MAC_0_87, output_MAC_0_88, output_MAC_0_89, 
		output_MAC_0_90, output_MAC_0_91, output_MAC_0_92, output_MAC_0_93, output_MAC_0_94, output_MAC_0_95, output_MAC_0_96, output_MAC_0_97, output_MAC_0_98, output_MAC_0_99, 
		output_MAC_0_100, output_MAC_0_101, output_MAC_0_102, output_MAC_0_103, output_MAC_0_104, output_MAC_0_105, output_MAC_0_106, output_MAC_0_107, output_MAC_0_108, output_MAC_0_109, 
		output_MAC_0_110, output_MAC_0_111, output_MAC_0_112, output_MAC_0_113, output_MAC_0_114, output_MAC_0_115, output_MAC_0_116, output_MAC_0_117, output_MAC_0_118, output_MAC_0_119, 
		output_MAC_0_120, output_MAC_0_121, output_MAC_0_122, output_MAC_0_123, output_MAC_0_124, output_MAC_0_125, output_MAC_0_126, output_MAC_0_127, output_MAC_0_128, output_MAC_0_129, 
		output_MAC_0_130, output_MAC_0_131, output_MAC_0_132, output_MAC_0_133, output_MAC_0_134, output_MAC_0_135, output_MAC_0_136, output_MAC_0_137, output_MAC_0_138, output_MAC_0_139, 
		output_MAC_0_140, output_MAC_0_141, output_MAC_0_142, output_MAC_0_143, output_MAC_0_144, output_MAC_0_145, output_MAC_0_146, output_MAC_0_147, output_MAC_0_148, output_MAC_0_149, 
		output_MAC_0_150, output_MAC_0_151, output_MAC_0_152, output_MAC_0_153, output_MAC_0_154, output_MAC_0_155, output_MAC_0_156, output_MAC_0_157, output_MAC_0_158, output_MAC_0_159, 
		output_MAC_0_160, output_MAC_0_161, output_MAC_0_162, output_MAC_0_163, output_MAC_0_164, output_MAC_0_165, output_MAC_0_166, output_MAC_0_167, output_MAC_0_168, output_MAC_0_169, 
		output_MAC_0_170, output_MAC_0_171, output_MAC_0_172, output_MAC_0_173, output_MAC_0_174, output_MAC_0_175, output_MAC_0_176, output_MAC_0_177, output_MAC_0_178, output_MAC_0_179, 
		output_MAC_0_180, output_MAC_0_181, output_MAC_0_182, output_MAC_0_183, output_MAC_0_184, output_MAC_0_185, output_MAC_0_186, output_MAC_0_187, output_MAC_0_188, output_MAC_0_189, 
		output_MAC_0_190, output_MAC_0_191, output_MAC_0_192, output_MAC_0_193, output_MAC_0_194, output_MAC_0_195, output_MAC_0_196, output_MAC_0_197, output_MAC_0_198, output_MAC_0_199, 
		output_MAC_0_200, output_MAC_0_201, output_MAC_0_202, output_MAC_0_203, output_MAC_0_204, output_MAC_0_205, output_MAC_0_206, output_MAC_0_207, output_MAC_0_208, output_MAC_0_209, 
		output_MAC_0_210, output_MAC_0_211, output_MAC_0_212, output_MAC_0_213, output_MAC_0_214, output_MAC_0_215, output_MAC_0_216, output_MAC_0_217, output_MAC_0_218, output_MAC_0_219, 
		output_MAC_0_220, output_MAC_0_221, output_MAC_0_222, output_MAC_0_223, output_MAC_0_224, output_MAC_0_225, output_MAC_0_226, output_MAC_0_227, output_MAC_0_228, output_MAC_0_229, 
		output_MAC_0_230, output_MAC_0_231, output_MAC_0_232, output_MAC_0_233, output_MAC_0_234, output_MAC_0_235, output_MAC_0_236, output_MAC_0_237, output_MAC_0_238, output_MAC_0_239, 
		output_MAC_0_240, output_MAC_0_241, output_MAC_0_242, output_MAC_0_243, output_MAC_0_244, output_MAC_0_245, output_MAC_0_246, output_MAC_0_247, output_MAC_0_248, output_MAC_0_249, 
		output_MAC_0_250, output_MAC_0_251, output_MAC_0_252, output_MAC_0_253, output_MAC_0_254, output_MAC_0_255, output_MAC_0_256, output_MAC_0_257, output_MAC_0_258, output_MAC_0_259, 
		output_MAC_0_260, output_MAC_0_261, output_MAC_0_262, output_MAC_0_263, output_MAC_0_264, output_MAC_0_265, output_MAC_0_266, output_MAC_0_267, output_MAC_0_268, output_MAC_0_269, 
		output_MAC_0_270, output_MAC_0_271, output_MAC_0_272, output_MAC_0_273, output_MAC_0_274, output_MAC_0_275, output_MAC_0_276, output_MAC_0_277, output_MAC_0_278, output_MAC_0_279, 
		output_MAC_0_280, output_MAC_0_281, output_MAC_0_282, output_MAC_0_283, output_MAC_0_284, output_MAC_0_285, output_MAC_0_286, output_MAC_0_287, output_MAC_0_288, output_MAC_0_289, 
		output_MAC_0_290, output_MAC_0_291, output_MAC_0_292, output_MAC_0_293, output_MAC_0_294, output_MAC_0_295, output_MAC_0_296, output_MAC_0_297, output_MAC_0_298, output_MAC_0_299, 
		output_MAC_0_300, output_MAC_0_301, output_MAC_0_302, output_MAC_0_303, output_MAC_0_304, output_MAC_0_305, output_MAC_0_306, output_MAC_0_307, output_MAC_0_308, output_MAC_0_309, 
		output_MAC_0_310, output_MAC_0_311, output_MAC_0_312, output_MAC_0_313, output_MAC_0_314, output_MAC_0_315, output_MAC_0_316, output_MAC_0_317, output_MAC_0_318, output_MAC_0_319, 
		output_MAC_0_320, output_MAC_0_321, output_MAC_0_322, output_MAC_0_323, output_MAC_0_324, output_MAC_0_325, output_MAC_0_326, output_MAC_0_327, output_MAC_0_328, output_MAC_0_329, 
		output_MAC_0_330, output_MAC_0_331, output_MAC_0_332, output_MAC_0_333, output_MAC_0_334, output_MAC_0_335, output_MAC_0_336, output_MAC_0_337, output_MAC_0_338, output_MAC_0_339, 
		output_MAC_0_340, output_MAC_0_341, output_MAC_0_342, output_MAC_0_343, output_MAC_0_344, output_MAC_0_345, output_MAC_0_346, output_MAC_0_347, output_MAC_0_348, output_MAC_0_349, 
		output_MAC_0_350, output_MAC_0_351, output_MAC_0_352, output_MAC_0_353, output_MAC_0_354, output_MAC_0_355, output_MAC_0_356, output_MAC_0_357, output_MAC_0_358, output_MAC_0_359, 
		output_MAC_0_360, output_MAC_0_361, output_MAC_0_362, output_MAC_0_363, output_MAC_0_364, output_MAC_0_365, output_MAC_0_366, output_MAC_0_367, output_MAC_0_368, output_MAC_0_369, 
		output_MAC_0_370, output_MAC_0_371, output_MAC_0_372, output_MAC_0_373, output_MAC_0_374, output_MAC_0_375, output_MAC_0_376, output_MAC_0_377, output_MAC_0_378, output_MAC_0_379, 
		output_MAC_0_380, output_MAC_0_381, output_MAC_0_382, output_MAC_0_383, output_MAC_0_384, output_MAC_0_385, output_MAC_0_386, output_MAC_0_387, output_MAC_0_388, output_MAC_0_389, 
		output_MAC_0_390, output_MAC_0_391, output_MAC_0_392, output_MAC_0_393, output_MAC_0_394, output_MAC_0_395, output_MAC_0_396, output_MAC_0_397, output_MAC_0_398, output_MAC_0_399, 
		output_MAC_0_400, output_MAC_0_401, output_MAC_0_402, output_MAC_0_403, output_MAC_0_404, output_MAC_0_405, output_MAC_0_406, output_MAC_0_407, output_MAC_0_408, output_MAC_0_409, 
		output_MAC_0_410, output_MAC_0_411, output_MAC_0_412, output_MAC_0_413, output_MAC_0_414, output_MAC_0_415, output_MAC_0_416, output_MAC_0_417, output_MAC_0_418, output_MAC_0_419, 
		output_MAC_0_420, output_MAC_0_421, output_MAC_0_422, output_MAC_0_423, output_MAC_0_424, output_MAC_0_425, output_MAC_0_426, output_MAC_0_427, output_MAC_0_428, output_MAC_0_429, 
		output_MAC_0_430, output_MAC_0_431, output_MAC_0_432, output_MAC_0_433, output_MAC_0_434, output_MAC_0_435, output_MAC_0_436, output_MAC_0_437, output_MAC_0_438, output_MAC_0_439, 
		output_MAC_0_440, output_MAC_0_441, output_MAC_0_442, output_MAC_0_443, output_MAC_0_444, output_MAC_0_445, output_MAC_0_446, output_MAC_0_447, output_MAC_0_448, output_MAC_0_449, 
		output_MAC_0_450, output_MAC_0_451, output_MAC_0_452, output_MAC_0_453, output_MAC_0_454, output_MAC_0_455, output_MAC_0_456, output_MAC_0_457, output_MAC_0_458, output_MAC_0_459, 
		output_MAC_0_460, output_MAC_0_461, output_MAC_0_462, output_MAC_0_463, output_MAC_0_464, output_MAC_0_465, output_MAC_0_466, output_MAC_0_467, output_MAC_0_468, output_MAC_0_469, 
		output_MAC_0_470, output_MAC_0_471, output_MAC_0_472, output_MAC_0_473, output_MAC_0_474, output_MAC_0_475, output_MAC_0_476, output_MAC_0_477, output_MAC_0_478, output_MAC_0_479, 
		output_MAC_0_480, output_MAC_0_481, output_MAC_0_482, output_MAC_0_483, output_MAC_0_484, output_MAC_0_485, output_MAC_0_486, output_MAC_0_487, output_MAC_0_488, output_MAC_0_489, 
		output_MAC_0_490, output_MAC_0_491, output_MAC_0_492, output_MAC_0_493, output_MAC_0_494, output_MAC_0_495, output_MAC_0_496, output_MAC_0_497, output_MAC_0_498, output_MAC_0_499, 
		output_MAC_0_500, output_MAC_0_501, output_MAC_0_502, output_MAC_0_503, output_MAC_0_504, output_MAC_0_505, output_MAC_0_506, output_MAC_0_507, output_MAC_0_508, output_MAC_0_509, 
		output_MAC_0_510, output_MAC_0_511, output_MAC_0_512, output_MAC_0_513, output_MAC_0_514, output_MAC_0_515, output_MAC_0_516, output_MAC_0_517, output_MAC_0_518, output_MAC_0_519, 
		output_MAC_0_520, output_MAC_0_521, output_MAC_0_522, output_MAC_0_523, output_MAC_0_524, output_MAC_0_525, output_MAC_0_526, output_MAC_0_527, output_MAC_0_528, output_MAC_0_529, 
		output_MAC_0_530, output_MAC_0_531, output_MAC_0_532, output_MAC_0_533, output_MAC_0_534, output_MAC_0_535, output_MAC_0_536, output_MAC_0_537, output_MAC_0_538, output_MAC_0_539, 
		output_MAC_0_540, output_MAC_0_541, output_MAC_0_542, output_MAC_0_543, output_MAC_0_544, output_MAC_0_545, output_MAC_0_546, output_MAC_0_547, output_MAC_0_548, output_MAC_0_549, 
		output_MAC_0_550, output_MAC_0_551, output_MAC_0_552, output_MAC_0_553, output_MAC_0_554, output_MAC_0_555, output_MAC_0_556, output_MAC_0_557, output_MAC_0_558, output_MAC_0_559, 
		output_MAC_0_560, output_MAC_0_561, output_MAC_0_562, output_MAC_0_563, output_MAC_0_564, output_MAC_0_565, output_MAC_0_566, output_MAC_0_567, output_MAC_0_568, output_MAC_0_569, 
		output_MAC_0_570, output_MAC_0_571, output_MAC_0_572, output_MAC_0_573, output_MAC_0_574, output_MAC_0_575, output_MAC_0_576, output_MAC_0_577, output_MAC_0_578, output_MAC_0_579, 
		output_MAC_0_580, output_MAC_0_581, output_MAC_0_582, output_MAC_0_583, output_MAC_0_584, output_MAC_0_585, output_MAC_0_586, output_MAC_0_587, output_MAC_0_588, output_MAC_0_589, 
		output_MAC_0_590, output_MAC_0_591, output_MAC_0_592, output_MAC_0_593, output_MAC_0_594, output_MAC_0_595, output_MAC_0_596, output_MAC_0_597, output_MAC_0_598, output_MAC_0_599, 
		output_MAC_0_600, output_MAC_0_601, output_MAC_0_602, output_MAC_0_603, output_MAC_0_604, output_MAC_0_605, output_MAC_0_606, output_MAC_0_607, output_MAC_0_608, output_MAC_0_609, 
		output_MAC_0_610, output_MAC_0_611, output_MAC_0_612, output_MAC_0_613, output_MAC_0_614, output_MAC_0_615, output_MAC_0_616, output_MAC_0_617, output_MAC_0_618, output_MAC_0_619, 
		output_MAC_0_620, output_MAC_0_621, output_MAC_0_622, output_MAC_0_623, output_MAC_0_624, output_MAC_0_625, output_MAC_0_626, output_MAC_0_627, output_MAC_0_628, output_MAC_0_629, 
		output_MAC_0_630, output_MAC_0_631, output_MAC_0_632, output_MAC_0_633, output_MAC_0_634, output_MAC_0_635, output_MAC_0_636, output_MAC_0_637, output_MAC_0_638, output_MAC_0_639, 
		output_MAC_0_640, output_MAC_0_641, output_MAC_0_642, output_MAC_0_643, output_MAC_0_644, output_MAC_0_645, output_MAC_0_646, output_MAC_0_647, output_MAC_0_648, output_MAC_0_649, 
		output_MAC_0_650, output_MAC_0_651, output_MAC_0_652, output_MAC_0_653, output_MAC_0_654, output_MAC_0_655, output_MAC_0_656, output_MAC_0_657, output_MAC_0_658, output_MAC_0_659, 
		output_MAC_0_660, output_MAC_0_661, output_MAC_0_662, output_MAC_0_663, output_MAC_0_664, output_MAC_0_665, output_MAC_0_666, output_MAC_0_667, output_MAC_0_668, output_MAC_0_669, 
		output_MAC_0_670, output_MAC_0_671, output_MAC_0_672, output_MAC_0_673, output_MAC_0_674, output_MAC_0_675, output_MAC_0_676, output_MAC_0_677, output_MAC_0_678, output_MAC_0_679, 
		output_MAC_0_680, output_MAC_0_681, output_MAC_0_682, output_MAC_0_683, output_MAC_0_684, output_MAC_0_685, output_MAC_0_686, output_MAC_0_687, output_MAC_0_688, output_MAC_0_689, 
		output_MAC_0_690, output_MAC_0_691, output_MAC_0_692, output_MAC_0_693, output_MAC_0_694, output_MAC_0_695, output_MAC_0_696, output_MAC_0_697, output_MAC_0_698, output_MAC_0_699, 
		output_MAC_0_700, output_MAC_0_701, output_MAC_0_702, output_MAC_0_703, output_MAC_0_704, output_MAC_0_705, output_MAC_0_706, output_MAC_0_707, output_MAC_0_708, output_MAC_0_709, 
		output_MAC_0_710, output_MAC_0_711, output_MAC_0_712, output_MAC_0_713, output_MAC_0_714, output_MAC_0_715, output_MAC_0_716, output_MAC_0_717, output_MAC_0_718, output_MAC_0_719, 
		output_MAC_0_720, output_MAC_0_721, output_MAC_0_722, output_MAC_0_723, output_MAC_0_724, output_MAC_0_725, output_MAC_0_726, output_MAC_0_727, output_MAC_0_728, output_MAC_0_729, 
		output_MAC_0_730, output_MAC_0_731, output_MAC_0_732, output_MAC_0_733, output_MAC_0_734, output_MAC_0_735, output_MAC_0_736, output_MAC_0_737, output_MAC_0_738, output_MAC_0_739, 
		output_MAC_0_740, output_MAC_0_741, output_MAC_0_742, output_MAC_0_743, output_MAC_0_744, output_MAC_0_745, output_MAC_0_746, output_MAC_0_747, output_MAC_0_748, output_MAC_0_749, 
		output_MAC_0_750, output_MAC_0_751, output_MAC_0_752, output_MAC_0_753, output_MAC_0_754, output_MAC_0_755, output_MAC_0_756, output_MAC_0_757, output_MAC_0_758, output_MAC_0_759, 
		output_MAC_0_760, output_MAC_0_761, output_MAC_0_762, output_MAC_0_763, output_MAC_0_764, output_MAC_0_765, output_MAC_0_766, output_MAC_0_767: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_1_0, output_MAC_1_1, output_MAC_1_2, output_MAC_1_3, output_MAC_1_4, output_MAC_1_5, output_MAC_1_6, output_MAC_1_7, output_MAC_1_8, output_MAC_1_9, 
		output_MAC_1_10, output_MAC_1_11, output_MAC_1_12, output_MAC_1_13, output_MAC_1_14, output_MAC_1_15, output_MAC_1_16, output_MAC_1_17, output_MAC_1_18, output_MAC_1_19, 
		output_MAC_1_20, output_MAC_1_21, output_MAC_1_22, output_MAC_1_23, output_MAC_1_24, output_MAC_1_25, output_MAC_1_26, output_MAC_1_27, output_MAC_1_28, output_MAC_1_29, 
		output_MAC_1_30, output_MAC_1_31, output_MAC_1_32, output_MAC_1_33, output_MAC_1_34, output_MAC_1_35, output_MAC_1_36, output_MAC_1_37, output_MAC_1_38, output_MAC_1_39, 
		output_MAC_1_40, output_MAC_1_41, output_MAC_1_42, output_MAC_1_43, output_MAC_1_44, output_MAC_1_45, output_MAC_1_46, output_MAC_1_47, output_MAC_1_48, output_MAC_1_49, 
		output_MAC_1_50, output_MAC_1_51, output_MAC_1_52, output_MAC_1_53, output_MAC_1_54, output_MAC_1_55, output_MAC_1_56, output_MAC_1_57, output_MAC_1_58, output_MAC_1_59, 
		output_MAC_1_60, output_MAC_1_61, output_MAC_1_62, output_MAC_1_63, output_MAC_1_64, output_MAC_1_65, output_MAC_1_66, output_MAC_1_67, output_MAC_1_68, output_MAC_1_69, 
		output_MAC_1_70, output_MAC_1_71, output_MAC_1_72, output_MAC_1_73, output_MAC_1_74, output_MAC_1_75, output_MAC_1_76, output_MAC_1_77, output_MAC_1_78, output_MAC_1_79, 
		output_MAC_1_80, output_MAC_1_81, output_MAC_1_82, output_MAC_1_83, output_MAC_1_84, output_MAC_1_85, output_MAC_1_86, output_MAC_1_87, output_MAC_1_88, output_MAC_1_89, 
		output_MAC_1_90, output_MAC_1_91, output_MAC_1_92, output_MAC_1_93, output_MAC_1_94, output_MAC_1_95, output_MAC_1_96, output_MAC_1_97, output_MAC_1_98, output_MAC_1_99, 
		output_MAC_1_100, output_MAC_1_101, output_MAC_1_102, output_MAC_1_103, output_MAC_1_104, output_MAC_1_105, output_MAC_1_106, output_MAC_1_107, output_MAC_1_108, output_MAC_1_109, 
		output_MAC_1_110, output_MAC_1_111, output_MAC_1_112, output_MAC_1_113, output_MAC_1_114, output_MAC_1_115, output_MAC_1_116, output_MAC_1_117, output_MAC_1_118, output_MAC_1_119, 
		output_MAC_1_120, output_MAC_1_121, output_MAC_1_122, output_MAC_1_123, output_MAC_1_124, output_MAC_1_125, output_MAC_1_126, output_MAC_1_127, output_MAC_1_128, output_MAC_1_129, 
		output_MAC_1_130, output_MAC_1_131, output_MAC_1_132, output_MAC_1_133, output_MAC_1_134, output_MAC_1_135, output_MAC_1_136, output_MAC_1_137, output_MAC_1_138, output_MAC_1_139, 
		output_MAC_1_140, output_MAC_1_141, output_MAC_1_142, output_MAC_1_143, output_MAC_1_144, output_MAC_1_145, output_MAC_1_146, output_MAC_1_147, output_MAC_1_148, output_MAC_1_149, 
		output_MAC_1_150, output_MAC_1_151, output_MAC_1_152, output_MAC_1_153, output_MAC_1_154, output_MAC_1_155, output_MAC_1_156, output_MAC_1_157, output_MAC_1_158, output_MAC_1_159, 
		output_MAC_1_160, output_MAC_1_161, output_MAC_1_162, output_MAC_1_163, output_MAC_1_164, output_MAC_1_165, output_MAC_1_166, output_MAC_1_167, output_MAC_1_168, output_MAC_1_169, 
		output_MAC_1_170, output_MAC_1_171, output_MAC_1_172, output_MAC_1_173, output_MAC_1_174, output_MAC_1_175, output_MAC_1_176, output_MAC_1_177, output_MAC_1_178, output_MAC_1_179, 
		output_MAC_1_180, output_MAC_1_181, output_MAC_1_182, output_MAC_1_183, output_MAC_1_184, output_MAC_1_185, output_MAC_1_186, output_MAC_1_187, output_MAC_1_188, output_MAC_1_189, 
		output_MAC_1_190, output_MAC_1_191, output_MAC_1_192, output_MAC_1_193, output_MAC_1_194, output_MAC_1_195, output_MAC_1_196, output_MAC_1_197, output_MAC_1_198, output_MAC_1_199, 
		output_MAC_1_200, output_MAC_1_201, output_MAC_1_202, output_MAC_1_203, output_MAC_1_204, output_MAC_1_205, output_MAC_1_206, output_MAC_1_207, output_MAC_1_208, output_MAC_1_209, 
		output_MAC_1_210, output_MAC_1_211, output_MAC_1_212, output_MAC_1_213, output_MAC_1_214, output_MAC_1_215, output_MAC_1_216, output_MAC_1_217, output_MAC_1_218, output_MAC_1_219, 
		output_MAC_1_220, output_MAC_1_221, output_MAC_1_222, output_MAC_1_223, output_MAC_1_224, output_MAC_1_225, output_MAC_1_226, output_MAC_1_227, output_MAC_1_228, output_MAC_1_229, 
		output_MAC_1_230, output_MAC_1_231, output_MAC_1_232, output_MAC_1_233, output_MAC_1_234, output_MAC_1_235, output_MAC_1_236, output_MAC_1_237, output_MAC_1_238, output_MAC_1_239, 
		output_MAC_1_240, output_MAC_1_241, output_MAC_1_242, output_MAC_1_243, output_MAC_1_244, output_MAC_1_245, output_MAC_1_246, output_MAC_1_247, output_MAC_1_248, output_MAC_1_249, 
		output_MAC_1_250, output_MAC_1_251, output_MAC_1_252, output_MAC_1_253, output_MAC_1_254, output_MAC_1_255, output_MAC_1_256, output_MAC_1_257, output_MAC_1_258, output_MAC_1_259, 
		output_MAC_1_260, output_MAC_1_261, output_MAC_1_262, output_MAC_1_263, output_MAC_1_264, output_MAC_1_265, output_MAC_1_266, output_MAC_1_267, output_MAC_1_268, output_MAC_1_269, 
		output_MAC_1_270, output_MAC_1_271, output_MAC_1_272, output_MAC_1_273, output_MAC_1_274, output_MAC_1_275, output_MAC_1_276, output_MAC_1_277, output_MAC_1_278, output_MAC_1_279, 
		output_MAC_1_280, output_MAC_1_281, output_MAC_1_282, output_MAC_1_283, output_MAC_1_284, output_MAC_1_285, output_MAC_1_286, output_MAC_1_287, output_MAC_1_288, output_MAC_1_289, 
		output_MAC_1_290, output_MAC_1_291, output_MAC_1_292, output_MAC_1_293, output_MAC_1_294, output_MAC_1_295, output_MAC_1_296, output_MAC_1_297, output_MAC_1_298, output_MAC_1_299, 
		output_MAC_1_300, output_MAC_1_301, output_MAC_1_302, output_MAC_1_303, output_MAC_1_304, output_MAC_1_305, output_MAC_1_306, output_MAC_1_307, output_MAC_1_308, output_MAC_1_309, 
		output_MAC_1_310, output_MAC_1_311, output_MAC_1_312, output_MAC_1_313, output_MAC_1_314, output_MAC_1_315, output_MAC_1_316, output_MAC_1_317, output_MAC_1_318, output_MAC_1_319, 
		output_MAC_1_320, output_MAC_1_321, output_MAC_1_322, output_MAC_1_323, output_MAC_1_324, output_MAC_1_325, output_MAC_1_326, output_MAC_1_327, output_MAC_1_328, output_MAC_1_329, 
		output_MAC_1_330, output_MAC_1_331, output_MAC_1_332, output_MAC_1_333, output_MAC_1_334, output_MAC_1_335, output_MAC_1_336, output_MAC_1_337, output_MAC_1_338, output_MAC_1_339, 
		output_MAC_1_340, output_MAC_1_341, output_MAC_1_342, output_MAC_1_343, output_MAC_1_344, output_MAC_1_345, output_MAC_1_346, output_MAC_1_347, output_MAC_1_348, output_MAC_1_349, 
		output_MAC_1_350, output_MAC_1_351, output_MAC_1_352, output_MAC_1_353, output_MAC_1_354, output_MAC_1_355, output_MAC_1_356, output_MAC_1_357, output_MAC_1_358, output_MAC_1_359, 
		output_MAC_1_360, output_MAC_1_361, output_MAC_1_362, output_MAC_1_363, output_MAC_1_364, output_MAC_1_365, output_MAC_1_366, output_MAC_1_367, output_MAC_1_368, output_MAC_1_369, 
		output_MAC_1_370, output_MAC_1_371, output_MAC_1_372, output_MAC_1_373, output_MAC_1_374, output_MAC_1_375, output_MAC_1_376, output_MAC_1_377, output_MAC_1_378, output_MAC_1_379, 
		output_MAC_1_380, output_MAC_1_381, output_MAC_1_382, output_MAC_1_383, output_MAC_1_384, output_MAC_1_385, output_MAC_1_386, output_MAC_1_387, output_MAC_1_388, output_MAC_1_389, 
		output_MAC_1_390, output_MAC_1_391, output_MAC_1_392, output_MAC_1_393, output_MAC_1_394, output_MAC_1_395, output_MAC_1_396, output_MAC_1_397, output_MAC_1_398, output_MAC_1_399, 
		output_MAC_1_400, output_MAC_1_401, output_MAC_1_402, output_MAC_1_403, output_MAC_1_404, output_MAC_1_405, output_MAC_1_406, output_MAC_1_407, output_MAC_1_408, output_MAC_1_409, 
		output_MAC_1_410, output_MAC_1_411, output_MAC_1_412, output_MAC_1_413, output_MAC_1_414, output_MAC_1_415, output_MAC_1_416, output_MAC_1_417, output_MAC_1_418, output_MAC_1_419, 
		output_MAC_1_420, output_MAC_1_421, output_MAC_1_422, output_MAC_1_423, output_MAC_1_424, output_MAC_1_425, output_MAC_1_426, output_MAC_1_427, output_MAC_1_428, output_MAC_1_429, 
		output_MAC_1_430, output_MAC_1_431, output_MAC_1_432, output_MAC_1_433, output_MAC_1_434, output_MAC_1_435, output_MAC_1_436, output_MAC_1_437, output_MAC_1_438, output_MAC_1_439, 
		output_MAC_1_440, output_MAC_1_441, output_MAC_1_442, output_MAC_1_443, output_MAC_1_444, output_MAC_1_445, output_MAC_1_446, output_MAC_1_447, output_MAC_1_448, output_MAC_1_449, 
		output_MAC_1_450, output_MAC_1_451, output_MAC_1_452, output_MAC_1_453, output_MAC_1_454, output_MAC_1_455, output_MAC_1_456, output_MAC_1_457, output_MAC_1_458, output_MAC_1_459, 
		output_MAC_1_460, output_MAC_1_461, output_MAC_1_462, output_MAC_1_463, output_MAC_1_464, output_MAC_1_465, output_MAC_1_466, output_MAC_1_467, output_MAC_1_468, output_MAC_1_469, 
		output_MAC_1_470, output_MAC_1_471, output_MAC_1_472, output_MAC_1_473, output_MAC_1_474, output_MAC_1_475, output_MAC_1_476, output_MAC_1_477, output_MAC_1_478, output_MAC_1_479, 
		output_MAC_1_480, output_MAC_1_481, output_MAC_1_482, output_MAC_1_483, output_MAC_1_484, output_MAC_1_485, output_MAC_1_486, output_MAC_1_487, output_MAC_1_488, output_MAC_1_489, 
		output_MAC_1_490, output_MAC_1_491, output_MAC_1_492, output_MAC_1_493, output_MAC_1_494, output_MAC_1_495, output_MAC_1_496, output_MAC_1_497, output_MAC_1_498, output_MAC_1_499, 
		output_MAC_1_500, output_MAC_1_501, output_MAC_1_502, output_MAC_1_503, output_MAC_1_504, output_MAC_1_505, output_MAC_1_506, output_MAC_1_507, output_MAC_1_508, output_MAC_1_509, 
		output_MAC_1_510, output_MAC_1_511, output_MAC_1_512, output_MAC_1_513, output_MAC_1_514, output_MAC_1_515, output_MAC_1_516, output_MAC_1_517, output_MAC_1_518, output_MAC_1_519, 
		output_MAC_1_520, output_MAC_1_521, output_MAC_1_522, output_MAC_1_523, output_MAC_1_524, output_MAC_1_525, output_MAC_1_526, output_MAC_1_527, output_MAC_1_528, output_MAC_1_529, 
		output_MAC_1_530, output_MAC_1_531, output_MAC_1_532, output_MAC_1_533, output_MAC_1_534, output_MAC_1_535, output_MAC_1_536, output_MAC_1_537, output_MAC_1_538, output_MAC_1_539, 
		output_MAC_1_540, output_MAC_1_541, output_MAC_1_542, output_MAC_1_543, output_MAC_1_544, output_MAC_1_545, output_MAC_1_546, output_MAC_1_547, output_MAC_1_548, output_MAC_1_549, 
		output_MAC_1_550, output_MAC_1_551, output_MAC_1_552, output_MAC_1_553, output_MAC_1_554, output_MAC_1_555, output_MAC_1_556, output_MAC_1_557, output_MAC_1_558, output_MAC_1_559, 
		output_MAC_1_560, output_MAC_1_561, output_MAC_1_562, output_MAC_1_563, output_MAC_1_564, output_MAC_1_565, output_MAC_1_566, output_MAC_1_567, output_MAC_1_568, output_MAC_1_569, 
		output_MAC_1_570, output_MAC_1_571, output_MAC_1_572, output_MAC_1_573, output_MAC_1_574, output_MAC_1_575, output_MAC_1_576, output_MAC_1_577, output_MAC_1_578, output_MAC_1_579, 
		output_MAC_1_580, output_MAC_1_581, output_MAC_1_582, output_MAC_1_583, output_MAC_1_584, output_MAC_1_585, output_MAC_1_586, output_MAC_1_587, output_MAC_1_588, output_MAC_1_589, 
		output_MAC_1_590, output_MAC_1_591, output_MAC_1_592, output_MAC_1_593, output_MAC_1_594, output_MAC_1_595, output_MAC_1_596, output_MAC_1_597, output_MAC_1_598, output_MAC_1_599, 
		output_MAC_1_600, output_MAC_1_601, output_MAC_1_602, output_MAC_1_603, output_MAC_1_604, output_MAC_1_605, output_MAC_1_606, output_MAC_1_607, output_MAC_1_608, output_MAC_1_609, 
		output_MAC_1_610, output_MAC_1_611, output_MAC_1_612, output_MAC_1_613, output_MAC_1_614, output_MAC_1_615, output_MAC_1_616, output_MAC_1_617, output_MAC_1_618, output_MAC_1_619, 
		output_MAC_1_620, output_MAC_1_621, output_MAC_1_622, output_MAC_1_623, output_MAC_1_624, output_MAC_1_625, output_MAC_1_626, output_MAC_1_627, output_MAC_1_628, output_MAC_1_629, 
		output_MAC_1_630, output_MAC_1_631, output_MAC_1_632, output_MAC_1_633, output_MAC_1_634, output_MAC_1_635, output_MAC_1_636, output_MAC_1_637, output_MAC_1_638, output_MAC_1_639, 
		output_MAC_1_640, output_MAC_1_641, output_MAC_1_642, output_MAC_1_643, output_MAC_1_644, output_MAC_1_645, output_MAC_1_646, output_MAC_1_647, output_MAC_1_648, output_MAC_1_649, 
		output_MAC_1_650, output_MAC_1_651, output_MAC_1_652, output_MAC_1_653, output_MAC_1_654, output_MAC_1_655, output_MAC_1_656, output_MAC_1_657, output_MAC_1_658, output_MAC_1_659, 
		output_MAC_1_660, output_MAC_1_661, output_MAC_1_662, output_MAC_1_663, output_MAC_1_664, output_MAC_1_665, output_MAC_1_666, output_MAC_1_667, output_MAC_1_668, output_MAC_1_669, 
		output_MAC_1_670, output_MAC_1_671, output_MAC_1_672, output_MAC_1_673, output_MAC_1_674, output_MAC_1_675, output_MAC_1_676, output_MAC_1_677, output_MAC_1_678, output_MAC_1_679, 
		output_MAC_1_680, output_MAC_1_681, output_MAC_1_682, output_MAC_1_683, output_MAC_1_684, output_MAC_1_685, output_MAC_1_686, output_MAC_1_687, output_MAC_1_688, output_MAC_1_689, 
		output_MAC_1_690, output_MAC_1_691, output_MAC_1_692, output_MAC_1_693, output_MAC_1_694, output_MAC_1_695, output_MAC_1_696, output_MAC_1_697, output_MAC_1_698, output_MAC_1_699, 
		output_MAC_1_700, output_MAC_1_701, output_MAC_1_702, output_MAC_1_703, output_MAC_1_704, output_MAC_1_705, output_MAC_1_706, output_MAC_1_707, output_MAC_1_708, output_MAC_1_709, 
		output_MAC_1_710, output_MAC_1_711, output_MAC_1_712, output_MAC_1_713, output_MAC_1_714, output_MAC_1_715, output_MAC_1_716, output_MAC_1_717, output_MAC_1_718, output_MAC_1_719, 
		output_MAC_1_720, output_MAC_1_721, output_MAC_1_722, output_MAC_1_723, output_MAC_1_724, output_MAC_1_725, output_MAC_1_726, output_MAC_1_727, output_MAC_1_728, output_MAC_1_729, 
		output_MAC_1_730, output_MAC_1_731, output_MAC_1_732, output_MAC_1_733, output_MAC_1_734, output_MAC_1_735, output_MAC_1_736, output_MAC_1_737, output_MAC_1_738, output_MAC_1_739, 
		output_MAC_1_740, output_MAC_1_741, output_MAC_1_742, output_MAC_1_743, output_MAC_1_744, output_MAC_1_745, output_MAC_1_746, output_MAC_1_747, output_MAC_1_748, output_MAC_1_749, 
		output_MAC_1_750, output_MAC_1_751, output_MAC_1_752, output_MAC_1_753, output_MAC_1_754, output_MAC_1_755, output_MAC_1_756, output_MAC_1_757, output_MAC_1_758, output_MAC_1_759, 
		output_MAC_1_760, output_MAC_1_761, output_MAC_1_762, output_MAC_1_763, output_MAC_1_764, output_MAC_1_765, output_MAC_1_766, output_MAC_1_767: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_2_0, output_MAC_2_1, output_MAC_2_2, output_MAC_2_3, output_MAC_2_4, output_MAC_2_5, output_MAC_2_6, output_MAC_2_7, output_MAC_2_8, output_MAC_2_9, 
		output_MAC_2_10, output_MAC_2_11, output_MAC_2_12, output_MAC_2_13, output_MAC_2_14, output_MAC_2_15, output_MAC_2_16, output_MAC_2_17, output_MAC_2_18, output_MAC_2_19, 
		output_MAC_2_20, output_MAC_2_21, output_MAC_2_22, output_MAC_2_23, output_MAC_2_24, output_MAC_2_25, output_MAC_2_26, output_MAC_2_27, output_MAC_2_28, output_MAC_2_29, 
		output_MAC_2_30, output_MAC_2_31, output_MAC_2_32, output_MAC_2_33, output_MAC_2_34, output_MAC_2_35, output_MAC_2_36, output_MAC_2_37, output_MAC_2_38, output_MAC_2_39, 
		output_MAC_2_40, output_MAC_2_41, output_MAC_2_42, output_MAC_2_43, output_MAC_2_44, output_MAC_2_45, output_MAC_2_46, output_MAC_2_47, output_MAC_2_48, output_MAC_2_49, 
		output_MAC_2_50, output_MAC_2_51, output_MAC_2_52, output_MAC_2_53, output_MAC_2_54, output_MAC_2_55, output_MAC_2_56, output_MAC_2_57, output_MAC_2_58, output_MAC_2_59, 
		output_MAC_2_60, output_MAC_2_61, output_MAC_2_62, output_MAC_2_63, output_MAC_2_64, output_MAC_2_65, output_MAC_2_66, output_MAC_2_67, output_MAC_2_68, output_MAC_2_69, 
		output_MAC_2_70, output_MAC_2_71, output_MAC_2_72, output_MAC_2_73, output_MAC_2_74, output_MAC_2_75, output_MAC_2_76, output_MAC_2_77, output_MAC_2_78, output_MAC_2_79, 
		output_MAC_2_80, output_MAC_2_81, output_MAC_2_82, output_MAC_2_83, output_MAC_2_84, output_MAC_2_85, output_MAC_2_86, output_MAC_2_87, output_MAC_2_88, output_MAC_2_89, 
		output_MAC_2_90, output_MAC_2_91, output_MAC_2_92, output_MAC_2_93, output_MAC_2_94, output_MAC_2_95, output_MAC_2_96, output_MAC_2_97, output_MAC_2_98, output_MAC_2_99, 
		output_MAC_2_100, output_MAC_2_101, output_MAC_2_102, output_MAC_2_103, output_MAC_2_104, output_MAC_2_105, output_MAC_2_106, output_MAC_2_107, output_MAC_2_108, output_MAC_2_109, 
		output_MAC_2_110, output_MAC_2_111, output_MAC_2_112, output_MAC_2_113, output_MAC_2_114, output_MAC_2_115, output_MAC_2_116, output_MAC_2_117, output_MAC_2_118, output_MAC_2_119, 
		output_MAC_2_120, output_MAC_2_121, output_MAC_2_122, output_MAC_2_123, output_MAC_2_124, output_MAC_2_125, output_MAC_2_126, output_MAC_2_127, output_MAC_2_128, output_MAC_2_129, 
		output_MAC_2_130, output_MAC_2_131, output_MAC_2_132, output_MAC_2_133, output_MAC_2_134, output_MAC_2_135, output_MAC_2_136, output_MAC_2_137, output_MAC_2_138, output_MAC_2_139, 
		output_MAC_2_140, output_MAC_2_141, output_MAC_2_142, output_MAC_2_143, output_MAC_2_144, output_MAC_2_145, output_MAC_2_146, output_MAC_2_147, output_MAC_2_148, output_MAC_2_149, 
		output_MAC_2_150, output_MAC_2_151, output_MAC_2_152, output_MAC_2_153, output_MAC_2_154, output_MAC_2_155, output_MAC_2_156, output_MAC_2_157, output_MAC_2_158, output_MAC_2_159, 
		output_MAC_2_160, output_MAC_2_161, output_MAC_2_162, output_MAC_2_163, output_MAC_2_164, output_MAC_2_165, output_MAC_2_166, output_MAC_2_167, output_MAC_2_168, output_MAC_2_169, 
		output_MAC_2_170, output_MAC_2_171, output_MAC_2_172, output_MAC_2_173, output_MAC_2_174, output_MAC_2_175, output_MAC_2_176, output_MAC_2_177, output_MAC_2_178, output_MAC_2_179, 
		output_MAC_2_180, output_MAC_2_181, output_MAC_2_182, output_MAC_2_183, output_MAC_2_184, output_MAC_2_185, output_MAC_2_186, output_MAC_2_187, output_MAC_2_188, output_MAC_2_189, 
		output_MAC_2_190, output_MAC_2_191, output_MAC_2_192, output_MAC_2_193, output_MAC_2_194, output_MAC_2_195, output_MAC_2_196, output_MAC_2_197, output_MAC_2_198, output_MAC_2_199, 
		output_MAC_2_200, output_MAC_2_201, output_MAC_2_202, output_MAC_2_203, output_MAC_2_204, output_MAC_2_205, output_MAC_2_206, output_MAC_2_207, output_MAC_2_208, output_MAC_2_209, 
		output_MAC_2_210, output_MAC_2_211, output_MAC_2_212, output_MAC_2_213, output_MAC_2_214, output_MAC_2_215, output_MAC_2_216, output_MAC_2_217, output_MAC_2_218, output_MAC_2_219, 
		output_MAC_2_220, output_MAC_2_221, output_MAC_2_222, output_MAC_2_223, output_MAC_2_224, output_MAC_2_225, output_MAC_2_226, output_MAC_2_227, output_MAC_2_228, output_MAC_2_229, 
		output_MAC_2_230, output_MAC_2_231, output_MAC_2_232, output_MAC_2_233, output_MAC_2_234, output_MAC_2_235, output_MAC_2_236, output_MAC_2_237, output_MAC_2_238, output_MAC_2_239, 
		output_MAC_2_240, output_MAC_2_241, output_MAC_2_242, output_MAC_2_243, output_MAC_2_244, output_MAC_2_245, output_MAC_2_246, output_MAC_2_247, output_MAC_2_248, output_MAC_2_249, 
		output_MAC_2_250, output_MAC_2_251, output_MAC_2_252, output_MAC_2_253, output_MAC_2_254, output_MAC_2_255, output_MAC_2_256, output_MAC_2_257, output_MAC_2_258, output_MAC_2_259, 
		output_MAC_2_260, output_MAC_2_261, output_MAC_2_262, output_MAC_2_263, output_MAC_2_264, output_MAC_2_265, output_MAC_2_266, output_MAC_2_267, output_MAC_2_268, output_MAC_2_269, 
		output_MAC_2_270, output_MAC_2_271, output_MAC_2_272, output_MAC_2_273, output_MAC_2_274, output_MAC_2_275, output_MAC_2_276, output_MAC_2_277, output_MAC_2_278, output_MAC_2_279, 
		output_MAC_2_280, output_MAC_2_281, output_MAC_2_282, output_MAC_2_283, output_MAC_2_284, output_MAC_2_285, output_MAC_2_286, output_MAC_2_287, output_MAC_2_288, output_MAC_2_289, 
		output_MAC_2_290, output_MAC_2_291, output_MAC_2_292, output_MAC_2_293, output_MAC_2_294, output_MAC_2_295, output_MAC_2_296, output_MAC_2_297, output_MAC_2_298, output_MAC_2_299, 
		output_MAC_2_300, output_MAC_2_301, output_MAC_2_302, output_MAC_2_303, output_MAC_2_304, output_MAC_2_305, output_MAC_2_306, output_MAC_2_307, output_MAC_2_308, output_MAC_2_309, 
		output_MAC_2_310, output_MAC_2_311, output_MAC_2_312, output_MAC_2_313, output_MAC_2_314, output_MAC_2_315, output_MAC_2_316, output_MAC_2_317, output_MAC_2_318, output_MAC_2_319, 
		output_MAC_2_320, output_MAC_2_321, output_MAC_2_322, output_MAC_2_323, output_MAC_2_324, output_MAC_2_325, output_MAC_2_326, output_MAC_2_327, output_MAC_2_328, output_MAC_2_329, 
		output_MAC_2_330, output_MAC_2_331, output_MAC_2_332, output_MAC_2_333, output_MAC_2_334, output_MAC_2_335, output_MAC_2_336, output_MAC_2_337, output_MAC_2_338, output_MAC_2_339, 
		output_MAC_2_340, output_MAC_2_341, output_MAC_2_342, output_MAC_2_343, output_MAC_2_344, output_MAC_2_345, output_MAC_2_346, output_MAC_2_347, output_MAC_2_348, output_MAC_2_349, 
		output_MAC_2_350, output_MAC_2_351, output_MAC_2_352, output_MAC_2_353, output_MAC_2_354, output_MAC_2_355, output_MAC_2_356, output_MAC_2_357, output_MAC_2_358, output_MAC_2_359, 
		output_MAC_2_360, output_MAC_2_361, output_MAC_2_362, output_MAC_2_363, output_MAC_2_364, output_MAC_2_365, output_MAC_2_366, output_MAC_2_367, output_MAC_2_368, output_MAC_2_369, 
		output_MAC_2_370, output_MAC_2_371, output_MAC_2_372, output_MAC_2_373, output_MAC_2_374, output_MAC_2_375, output_MAC_2_376, output_MAC_2_377, output_MAC_2_378, output_MAC_2_379, 
		output_MAC_2_380, output_MAC_2_381, output_MAC_2_382, output_MAC_2_383, output_MAC_2_384, output_MAC_2_385, output_MAC_2_386, output_MAC_2_387, output_MAC_2_388, output_MAC_2_389, 
		output_MAC_2_390, output_MAC_2_391, output_MAC_2_392, output_MAC_2_393, output_MAC_2_394, output_MAC_2_395, output_MAC_2_396, output_MAC_2_397, output_MAC_2_398, output_MAC_2_399, 
		output_MAC_2_400, output_MAC_2_401, output_MAC_2_402, output_MAC_2_403, output_MAC_2_404, output_MAC_2_405, output_MAC_2_406, output_MAC_2_407, output_MAC_2_408, output_MAC_2_409, 
		output_MAC_2_410, output_MAC_2_411, output_MAC_2_412, output_MAC_2_413, output_MAC_2_414, output_MAC_2_415, output_MAC_2_416, output_MAC_2_417, output_MAC_2_418, output_MAC_2_419, 
		output_MAC_2_420, output_MAC_2_421, output_MAC_2_422, output_MAC_2_423, output_MAC_2_424, output_MAC_2_425, output_MAC_2_426, output_MAC_2_427, output_MAC_2_428, output_MAC_2_429, 
		output_MAC_2_430, output_MAC_2_431, output_MAC_2_432, output_MAC_2_433, output_MAC_2_434, output_MAC_2_435, output_MAC_2_436, output_MAC_2_437, output_MAC_2_438, output_MAC_2_439, 
		output_MAC_2_440, output_MAC_2_441, output_MAC_2_442, output_MAC_2_443, output_MAC_2_444, output_MAC_2_445, output_MAC_2_446, output_MAC_2_447, output_MAC_2_448, output_MAC_2_449, 
		output_MAC_2_450, output_MAC_2_451, output_MAC_2_452, output_MAC_2_453, output_MAC_2_454, output_MAC_2_455, output_MAC_2_456, output_MAC_2_457, output_MAC_2_458, output_MAC_2_459, 
		output_MAC_2_460, output_MAC_2_461, output_MAC_2_462, output_MAC_2_463, output_MAC_2_464, output_MAC_2_465, output_MAC_2_466, output_MAC_2_467, output_MAC_2_468, output_MAC_2_469, 
		output_MAC_2_470, output_MAC_2_471, output_MAC_2_472, output_MAC_2_473, output_MAC_2_474, output_MAC_2_475, output_MAC_2_476, output_MAC_2_477, output_MAC_2_478, output_MAC_2_479, 
		output_MAC_2_480, output_MAC_2_481, output_MAC_2_482, output_MAC_2_483, output_MAC_2_484, output_MAC_2_485, output_MAC_2_486, output_MAC_2_487, output_MAC_2_488, output_MAC_2_489, 
		output_MAC_2_490, output_MAC_2_491, output_MAC_2_492, output_MAC_2_493, output_MAC_2_494, output_MAC_2_495, output_MAC_2_496, output_MAC_2_497, output_MAC_2_498, output_MAC_2_499, 
		output_MAC_2_500, output_MAC_2_501, output_MAC_2_502, output_MAC_2_503, output_MAC_2_504, output_MAC_2_505, output_MAC_2_506, output_MAC_2_507, output_MAC_2_508, output_MAC_2_509, 
		output_MAC_2_510, output_MAC_2_511, output_MAC_2_512, output_MAC_2_513, output_MAC_2_514, output_MAC_2_515, output_MAC_2_516, output_MAC_2_517, output_MAC_2_518, output_MAC_2_519, 
		output_MAC_2_520, output_MAC_2_521, output_MAC_2_522, output_MAC_2_523, output_MAC_2_524, output_MAC_2_525, output_MAC_2_526, output_MAC_2_527, output_MAC_2_528, output_MAC_2_529, 
		output_MAC_2_530, output_MAC_2_531, output_MAC_2_532, output_MAC_2_533, output_MAC_2_534, output_MAC_2_535, output_MAC_2_536, output_MAC_2_537, output_MAC_2_538, output_MAC_2_539, 
		output_MAC_2_540, output_MAC_2_541, output_MAC_2_542, output_MAC_2_543, output_MAC_2_544, output_MAC_2_545, output_MAC_2_546, output_MAC_2_547, output_MAC_2_548, output_MAC_2_549, 
		output_MAC_2_550, output_MAC_2_551, output_MAC_2_552, output_MAC_2_553, output_MAC_2_554, output_MAC_2_555, output_MAC_2_556, output_MAC_2_557, output_MAC_2_558, output_MAC_2_559, 
		output_MAC_2_560, output_MAC_2_561, output_MAC_2_562, output_MAC_2_563, output_MAC_2_564, output_MAC_2_565, output_MAC_2_566, output_MAC_2_567, output_MAC_2_568, output_MAC_2_569, 
		output_MAC_2_570, output_MAC_2_571, output_MAC_2_572, output_MAC_2_573, output_MAC_2_574, output_MAC_2_575, output_MAC_2_576, output_MAC_2_577, output_MAC_2_578, output_MAC_2_579, 
		output_MAC_2_580, output_MAC_2_581, output_MAC_2_582, output_MAC_2_583, output_MAC_2_584, output_MAC_2_585, output_MAC_2_586, output_MAC_2_587, output_MAC_2_588, output_MAC_2_589, 
		output_MAC_2_590, output_MAC_2_591, output_MAC_2_592, output_MAC_2_593, output_MAC_2_594, output_MAC_2_595, output_MAC_2_596, output_MAC_2_597, output_MAC_2_598, output_MAC_2_599, 
		output_MAC_2_600, output_MAC_2_601, output_MAC_2_602, output_MAC_2_603, output_MAC_2_604, output_MAC_2_605, output_MAC_2_606, output_MAC_2_607, output_MAC_2_608, output_MAC_2_609, 
		output_MAC_2_610, output_MAC_2_611, output_MAC_2_612, output_MAC_2_613, output_MAC_2_614, output_MAC_2_615, output_MAC_2_616, output_MAC_2_617, output_MAC_2_618, output_MAC_2_619, 
		output_MAC_2_620, output_MAC_2_621, output_MAC_2_622, output_MAC_2_623, output_MAC_2_624, output_MAC_2_625, output_MAC_2_626, output_MAC_2_627, output_MAC_2_628, output_MAC_2_629, 
		output_MAC_2_630, output_MAC_2_631, output_MAC_2_632, output_MAC_2_633, output_MAC_2_634, output_MAC_2_635, output_MAC_2_636, output_MAC_2_637, output_MAC_2_638, output_MAC_2_639, 
		output_MAC_2_640, output_MAC_2_641, output_MAC_2_642, output_MAC_2_643, output_MAC_2_644, output_MAC_2_645, output_MAC_2_646, output_MAC_2_647, output_MAC_2_648, output_MAC_2_649, 
		output_MAC_2_650, output_MAC_2_651, output_MAC_2_652, output_MAC_2_653, output_MAC_2_654, output_MAC_2_655, output_MAC_2_656, output_MAC_2_657, output_MAC_2_658, output_MAC_2_659, 
		output_MAC_2_660, output_MAC_2_661, output_MAC_2_662, output_MAC_2_663, output_MAC_2_664, output_MAC_2_665, output_MAC_2_666, output_MAC_2_667, output_MAC_2_668, output_MAC_2_669, 
		output_MAC_2_670, output_MAC_2_671, output_MAC_2_672, output_MAC_2_673, output_MAC_2_674, output_MAC_2_675, output_MAC_2_676, output_MAC_2_677, output_MAC_2_678, output_MAC_2_679, 
		output_MAC_2_680, output_MAC_2_681, output_MAC_2_682, output_MAC_2_683, output_MAC_2_684, output_MAC_2_685, output_MAC_2_686, output_MAC_2_687, output_MAC_2_688, output_MAC_2_689, 
		output_MAC_2_690, output_MAC_2_691, output_MAC_2_692, output_MAC_2_693, output_MAC_2_694, output_MAC_2_695, output_MAC_2_696, output_MAC_2_697, output_MAC_2_698, output_MAC_2_699, 
		output_MAC_2_700, output_MAC_2_701, output_MAC_2_702, output_MAC_2_703, output_MAC_2_704, output_MAC_2_705, output_MAC_2_706, output_MAC_2_707, output_MAC_2_708, output_MAC_2_709, 
		output_MAC_2_710, output_MAC_2_711, output_MAC_2_712, output_MAC_2_713, output_MAC_2_714, output_MAC_2_715, output_MAC_2_716, output_MAC_2_717, output_MAC_2_718, output_MAC_2_719, 
		output_MAC_2_720, output_MAC_2_721, output_MAC_2_722, output_MAC_2_723, output_MAC_2_724, output_MAC_2_725, output_MAC_2_726, output_MAC_2_727, output_MAC_2_728, output_MAC_2_729, 
		output_MAC_2_730, output_MAC_2_731, output_MAC_2_732, output_MAC_2_733, output_MAC_2_734, output_MAC_2_735, output_MAC_2_736, output_MAC_2_737, output_MAC_2_738, output_MAC_2_739, 
		output_MAC_2_740, output_MAC_2_741, output_MAC_2_742, output_MAC_2_743, output_MAC_2_744, output_MAC_2_745, output_MAC_2_746, output_MAC_2_747, output_MAC_2_748, output_MAC_2_749, 
		output_MAC_2_750, output_MAC_2_751, output_MAC_2_752, output_MAC_2_753, output_MAC_2_754, output_MAC_2_755, output_MAC_2_756, output_MAC_2_757, output_MAC_2_758, output_MAC_2_759, 
		output_MAC_2_760, output_MAC_2_761, output_MAC_2_762, output_MAC_2_763, output_MAC_2_764, output_MAC_2_765, output_MAC_2_766, output_MAC_2_767: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_3_0, output_MAC_3_1, output_MAC_3_2, output_MAC_3_3, output_MAC_3_4, output_MAC_3_5, output_MAC_3_6, output_MAC_3_7, output_MAC_3_8, output_MAC_3_9, 
		output_MAC_3_10, output_MAC_3_11, output_MAC_3_12, output_MAC_3_13, output_MAC_3_14, output_MAC_3_15, output_MAC_3_16, output_MAC_3_17, output_MAC_3_18, output_MAC_3_19, 
		output_MAC_3_20, output_MAC_3_21, output_MAC_3_22, output_MAC_3_23, output_MAC_3_24, output_MAC_3_25, output_MAC_3_26, output_MAC_3_27, output_MAC_3_28, output_MAC_3_29, 
		output_MAC_3_30, output_MAC_3_31, output_MAC_3_32, output_MAC_3_33, output_MAC_3_34, output_MAC_3_35, output_MAC_3_36, output_MAC_3_37, output_MAC_3_38, output_MAC_3_39, 
		output_MAC_3_40, output_MAC_3_41, output_MAC_3_42, output_MAC_3_43, output_MAC_3_44, output_MAC_3_45, output_MAC_3_46, output_MAC_3_47, output_MAC_3_48, output_MAC_3_49, 
		output_MAC_3_50, output_MAC_3_51, output_MAC_3_52, output_MAC_3_53, output_MAC_3_54, output_MAC_3_55, output_MAC_3_56, output_MAC_3_57, output_MAC_3_58, output_MAC_3_59, 
		output_MAC_3_60, output_MAC_3_61, output_MAC_3_62, output_MAC_3_63, output_MAC_3_64, output_MAC_3_65, output_MAC_3_66, output_MAC_3_67, output_MAC_3_68, output_MAC_3_69, 
		output_MAC_3_70, output_MAC_3_71, output_MAC_3_72, output_MAC_3_73, output_MAC_3_74, output_MAC_3_75, output_MAC_3_76, output_MAC_3_77, output_MAC_3_78, output_MAC_3_79, 
		output_MAC_3_80, output_MAC_3_81, output_MAC_3_82, output_MAC_3_83, output_MAC_3_84, output_MAC_3_85, output_MAC_3_86, output_MAC_3_87, output_MAC_3_88, output_MAC_3_89, 
		output_MAC_3_90, output_MAC_3_91, output_MAC_3_92, output_MAC_3_93, output_MAC_3_94, output_MAC_3_95, output_MAC_3_96, output_MAC_3_97, output_MAC_3_98, output_MAC_3_99, 
		output_MAC_3_100, output_MAC_3_101, output_MAC_3_102, output_MAC_3_103, output_MAC_3_104, output_MAC_3_105, output_MAC_3_106, output_MAC_3_107, output_MAC_3_108, output_MAC_3_109, 
		output_MAC_3_110, output_MAC_3_111, output_MAC_3_112, output_MAC_3_113, output_MAC_3_114, output_MAC_3_115, output_MAC_3_116, output_MAC_3_117, output_MAC_3_118, output_MAC_3_119, 
		output_MAC_3_120, output_MAC_3_121, output_MAC_3_122, output_MAC_3_123, output_MAC_3_124, output_MAC_3_125, output_MAC_3_126, output_MAC_3_127, output_MAC_3_128, output_MAC_3_129, 
		output_MAC_3_130, output_MAC_3_131, output_MAC_3_132, output_MAC_3_133, output_MAC_3_134, output_MAC_3_135, output_MAC_3_136, output_MAC_3_137, output_MAC_3_138, output_MAC_3_139, 
		output_MAC_3_140, output_MAC_3_141, output_MAC_3_142, output_MAC_3_143, output_MAC_3_144, output_MAC_3_145, output_MAC_3_146, output_MAC_3_147, output_MAC_3_148, output_MAC_3_149, 
		output_MAC_3_150, output_MAC_3_151, output_MAC_3_152, output_MAC_3_153, output_MAC_3_154, output_MAC_3_155, output_MAC_3_156, output_MAC_3_157, output_MAC_3_158, output_MAC_3_159, 
		output_MAC_3_160, output_MAC_3_161, output_MAC_3_162, output_MAC_3_163, output_MAC_3_164, output_MAC_3_165, output_MAC_3_166, output_MAC_3_167, output_MAC_3_168, output_MAC_3_169, 
		output_MAC_3_170, output_MAC_3_171, output_MAC_3_172, output_MAC_3_173, output_MAC_3_174, output_MAC_3_175, output_MAC_3_176, output_MAC_3_177, output_MAC_3_178, output_MAC_3_179, 
		output_MAC_3_180, output_MAC_3_181, output_MAC_3_182, output_MAC_3_183, output_MAC_3_184, output_MAC_3_185, output_MAC_3_186, output_MAC_3_187, output_MAC_3_188, output_MAC_3_189, 
		output_MAC_3_190, output_MAC_3_191, output_MAC_3_192, output_MAC_3_193, output_MAC_3_194, output_MAC_3_195, output_MAC_3_196, output_MAC_3_197, output_MAC_3_198, output_MAC_3_199, 
		output_MAC_3_200, output_MAC_3_201, output_MAC_3_202, output_MAC_3_203, output_MAC_3_204, output_MAC_3_205, output_MAC_3_206, output_MAC_3_207, output_MAC_3_208, output_MAC_3_209, 
		output_MAC_3_210, output_MAC_3_211, output_MAC_3_212, output_MAC_3_213, output_MAC_3_214, output_MAC_3_215, output_MAC_3_216, output_MAC_3_217, output_MAC_3_218, output_MAC_3_219, 
		output_MAC_3_220, output_MAC_3_221, output_MAC_3_222, output_MAC_3_223, output_MAC_3_224, output_MAC_3_225, output_MAC_3_226, output_MAC_3_227, output_MAC_3_228, output_MAC_3_229, 
		output_MAC_3_230, output_MAC_3_231, output_MAC_3_232, output_MAC_3_233, output_MAC_3_234, output_MAC_3_235, output_MAC_3_236, output_MAC_3_237, output_MAC_3_238, output_MAC_3_239, 
		output_MAC_3_240, output_MAC_3_241, output_MAC_3_242, output_MAC_3_243, output_MAC_3_244, output_MAC_3_245, output_MAC_3_246, output_MAC_3_247, output_MAC_3_248, output_MAC_3_249, 
		output_MAC_3_250, output_MAC_3_251, output_MAC_3_252, output_MAC_3_253, output_MAC_3_254, output_MAC_3_255, output_MAC_3_256, output_MAC_3_257, output_MAC_3_258, output_MAC_3_259, 
		output_MAC_3_260, output_MAC_3_261, output_MAC_3_262, output_MAC_3_263, output_MAC_3_264, output_MAC_3_265, output_MAC_3_266, output_MAC_3_267, output_MAC_3_268, output_MAC_3_269, 
		output_MAC_3_270, output_MAC_3_271, output_MAC_3_272, output_MAC_3_273, output_MAC_3_274, output_MAC_3_275, output_MAC_3_276, output_MAC_3_277, output_MAC_3_278, output_MAC_3_279, 
		output_MAC_3_280, output_MAC_3_281, output_MAC_3_282, output_MAC_3_283, output_MAC_3_284, output_MAC_3_285, output_MAC_3_286, output_MAC_3_287, output_MAC_3_288, output_MAC_3_289, 
		output_MAC_3_290, output_MAC_3_291, output_MAC_3_292, output_MAC_3_293, output_MAC_3_294, output_MAC_3_295, output_MAC_3_296, output_MAC_3_297, output_MAC_3_298, output_MAC_3_299, 
		output_MAC_3_300, output_MAC_3_301, output_MAC_3_302, output_MAC_3_303, output_MAC_3_304, output_MAC_3_305, output_MAC_3_306, output_MAC_3_307, output_MAC_3_308, output_MAC_3_309, 
		output_MAC_3_310, output_MAC_3_311, output_MAC_3_312, output_MAC_3_313, output_MAC_3_314, output_MAC_3_315, output_MAC_3_316, output_MAC_3_317, output_MAC_3_318, output_MAC_3_319, 
		output_MAC_3_320, output_MAC_3_321, output_MAC_3_322, output_MAC_3_323, output_MAC_3_324, output_MAC_3_325, output_MAC_3_326, output_MAC_3_327, output_MAC_3_328, output_MAC_3_329, 
		output_MAC_3_330, output_MAC_3_331, output_MAC_3_332, output_MAC_3_333, output_MAC_3_334, output_MAC_3_335, output_MAC_3_336, output_MAC_3_337, output_MAC_3_338, output_MAC_3_339, 
		output_MAC_3_340, output_MAC_3_341, output_MAC_3_342, output_MAC_3_343, output_MAC_3_344, output_MAC_3_345, output_MAC_3_346, output_MAC_3_347, output_MAC_3_348, output_MAC_3_349, 
		output_MAC_3_350, output_MAC_3_351, output_MAC_3_352, output_MAC_3_353, output_MAC_3_354, output_MAC_3_355, output_MAC_3_356, output_MAC_3_357, output_MAC_3_358, output_MAC_3_359, 
		output_MAC_3_360, output_MAC_3_361, output_MAC_3_362, output_MAC_3_363, output_MAC_3_364, output_MAC_3_365, output_MAC_3_366, output_MAC_3_367, output_MAC_3_368, output_MAC_3_369, 
		output_MAC_3_370, output_MAC_3_371, output_MAC_3_372, output_MAC_3_373, output_MAC_3_374, output_MAC_3_375, output_MAC_3_376, output_MAC_3_377, output_MAC_3_378, output_MAC_3_379, 
		output_MAC_3_380, output_MAC_3_381, output_MAC_3_382, output_MAC_3_383, output_MAC_3_384, output_MAC_3_385, output_MAC_3_386, output_MAC_3_387, output_MAC_3_388, output_MAC_3_389, 
		output_MAC_3_390, output_MAC_3_391, output_MAC_3_392, output_MAC_3_393, output_MAC_3_394, output_MAC_3_395, output_MAC_3_396, output_MAC_3_397, output_MAC_3_398, output_MAC_3_399, 
		output_MAC_3_400, output_MAC_3_401, output_MAC_3_402, output_MAC_3_403, output_MAC_3_404, output_MAC_3_405, output_MAC_3_406, output_MAC_3_407, output_MAC_3_408, output_MAC_3_409, 
		output_MAC_3_410, output_MAC_3_411, output_MAC_3_412, output_MAC_3_413, output_MAC_3_414, output_MAC_3_415, output_MAC_3_416, output_MAC_3_417, output_MAC_3_418, output_MAC_3_419, 
		output_MAC_3_420, output_MAC_3_421, output_MAC_3_422, output_MAC_3_423, output_MAC_3_424, output_MAC_3_425, output_MAC_3_426, output_MAC_3_427, output_MAC_3_428, output_MAC_3_429, 
		output_MAC_3_430, output_MAC_3_431, output_MAC_3_432, output_MAC_3_433, output_MAC_3_434, output_MAC_3_435, output_MAC_3_436, output_MAC_3_437, output_MAC_3_438, output_MAC_3_439, 
		output_MAC_3_440, output_MAC_3_441, output_MAC_3_442, output_MAC_3_443, output_MAC_3_444, output_MAC_3_445, output_MAC_3_446, output_MAC_3_447, output_MAC_3_448, output_MAC_3_449, 
		output_MAC_3_450, output_MAC_3_451, output_MAC_3_452, output_MAC_3_453, output_MAC_3_454, output_MAC_3_455, output_MAC_3_456, output_MAC_3_457, output_MAC_3_458, output_MAC_3_459, 
		output_MAC_3_460, output_MAC_3_461, output_MAC_3_462, output_MAC_3_463, output_MAC_3_464, output_MAC_3_465, output_MAC_3_466, output_MAC_3_467, output_MAC_3_468, output_MAC_3_469, 
		output_MAC_3_470, output_MAC_3_471, output_MAC_3_472, output_MAC_3_473, output_MAC_3_474, output_MAC_3_475, output_MAC_3_476, output_MAC_3_477, output_MAC_3_478, output_MAC_3_479, 
		output_MAC_3_480, output_MAC_3_481, output_MAC_3_482, output_MAC_3_483, output_MAC_3_484, output_MAC_3_485, output_MAC_3_486, output_MAC_3_487, output_MAC_3_488, output_MAC_3_489, 
		output_MAC_3_490, output_MAC_3_491, output_MAC_3_492, output_MAC_3_493, output_MAC_3_494, output_MAC_3_495, output_MAC_3_496, output_MAC_3_497, output_MAC_3_498, output_MAC_3_499, 
		output_MAC_3_500, output_MAC_3_501, output_MAC_3_502, output_MAC_3_503, output_MAC_3_504, output_MAC_3_505, output_MAC_3_506, output_MAC_3_507, output_MAC_3_508, output_MAC_3_509, 
		output_MAC_3_510, output_MAC_3_511, output_MAC_3_512, output_MAC_3_513, output_MAC_3_514, output_MAC_3_515, output_MAC_3_516, output_MAC_3_517, output_MAC_3_518, output_MAC_3_519, 
		output_MAC_3_520, output_MAC_3_521, output_MAC_3_522, output_MAC_3_523, output_MAC_3_524, output_MAC_3_525, output_MAC_3_526, output_MAC_3_527, output_MAC_3_528, output_MAC_3_529, 
		output_MAC_3_530, output_MAC_3_531, output_MAC_3_532, output_MAC_3_533, output_MAC_3_534, output_MAC_3_535, output_MAC_3_536, output_MAC_3_537, output_MAC_3_538, output_MAC_3_539, 
		output_MAC_3_540, output_MAC_3_541, output_MAC_3_542, output_MAC_3_543, output_MAC_3_544, output_MAC_3_545, output_MAC_3_546, output_MAC_3_547, output_MAC_3_548, output_MAC_3_549, 
		output_MAC_3_550, output_MAC_3_551, output_MAC_3_552, output_MAC_3_553, output_MAC_3_554, output_MAC_3_555, output_MAC_3_556, output_MAC_3_557, output_MAC_3_558, output_MAC_3_559, 
		output_MAC_3_560, output_MAC_3_561, output_MAC_3_562, output_MAC_3_563, output_MAC_3_564, output_MAC_3_565, output_MAC_3_566, output_MAC_3_567, output_MAC_3_568, output_MAC_3_569, 
		output_MAC_3_570, output_MAC_3_571, output_MAC_3_572, output_MAC_3_573, output_MAC_3_574, output_MAC_3_575, output_MAC_3_576, output_MAC_3_577, output_MAC_3_578, output_MAC_3_579, 
		output_MAC_3_580, output_MAC_3_581, output_MAC_3_582, output_MAC_3_583, output_MAC_3_584, output_MAC_3_585, output_MAC_3_586, output_MAC_3_587, output_MAC_3_588, output_MAC_3_589, 
		output_MAC_3_590, output_MAC_3_591, output_MAC_3_592, output_MAC_3_593, output_MAC_3_594, output_MAC_3_595, output_MAC_3_596, output_MAC_3_597, output_MAC_3_598, output_MAC_3_599, 
		output_MAC_3_600, output_MAC_3_601, output_MAC_3_602, output_MAC_3_603, output_MAC_3_604, output_MAC_3_605, output_MAC_3_606, output_MAC_3_607, output_MAC_3_608, output_MAC_3_609, 
		output_MAC_3_610, output_MAC_3_611, output_MAC_3_612, output_MAC_3_613, output_MAC_3_614, output_MAC_3_615, output_MAC_3_616, output_MAC_3_617, output_MAC_3_618, output_MAC_3_619, 
		output_MAC_3_620, output_MAC_3_621, output_MAC_3_622, output_MAC_3_623, output_MAC_3_624, output_MAC_3_625, output_MAC_3_626, output_MAC_3_627, output_MAC_3_628, output_MAC_3_629, 
		output_MAC_3_630, output_MAC_3_631, output_MAC_3_632, output_MAC_3_633, output_MAC_3_634, output_MAC_3_635, output_MAC_3_636, output_MAC_3_637, output_MAC_3_638, output_MAC_3_639, 
		output_MAC_3_640, output_MAC_3_641, output_MAC_3_642, output_MAC_3_643, output_MAC_3_644, output_MAC_3_645, output_MAC_3_646, output_MAC_3_647, output_MAC_3_648, output_MAC_3_649, 
		output_MAC_3_650, output_MAC_3_651, output_MAC_3_652, output_MAC_3_653, output_MAC_3_654, output_MAC_3_655, output_MAC_3_656, output_MAC_3_657, output_MAC_3_658, output_MAC_3_659, 
		output_MAC_3_660, output_MAC_3_661, output_MAC_3_662, output_MAC_3_663, output_MAC_3_664, output_MAC_3_665, output_MAC_3_666, output_MAC_3_667, output_MAC_3_668, output_MAC_3_669, 
		output_MAC_3_670, output_MAC_3_671, output_MAC_3_672, output_MAC_3_673, output_MAC_3_674, output_MAC_3_675, output_MAC_3_676, output_MAC_3_677, output_MAC_3_678, output_MAC_3_679, 
		output_MAC_3_680, output_MAC_3_681, output_MAC_3_682, output_MAC_3_683, output_MAC_3_684, output_MAC_3_685, output_MAC_3_686, output_MAC_3_687, output_MAC_3_688, output_MAC_3_689, 
		output_MAC_3_690, output_MAC_3_691, output_MAC_3_692, output_MAC_3_693, output_MAC_3_694, output_MAC_3_695, output_MAC_3_696, output_MAC_3_697, output_MAC_3_698, output_MAC_3_699, 
		output_MAC_3_700, output_MAC_3_701, output_MAC_3_702, output_MAC_3_703, output_MAC_3_704, output_MAC_3_705, output_MAC_3_706, output_MAC_3_707, output_MAC_3_708, output_MAC_3_709, 
		output_MAC_3_710, output_MAC_3_711, output_MAC_3_712, output_MAC_3_713, output_MAC_3_714, output_MAC_3_715, output_MAC_3_716, output_MAC_3_717, output_MAC_3_718, output_MAC_3_719, 
		output_MAC_3_720, output_MAC_3_721, output_MAC_3_722, output_MAC_3_723, output_MAC_3_724, output_MAC_3_725, output_MAC_3_726, output_MAC_3_727, output_MAC_3_728, output_MAC_3_729, 
		output_MAC_3_730, output_MAC_3_731, output_MAC_3_732, output_MAC_3_733, output_MAC_3_734, output_MAC_3_735, output_MAC_3_736, output_MAC_3_737, output_MAC_3_738, output_MAC_3_739, 
		output_MAC_3_740, output_MAC_3_741, output_MAC_3_742, output_MAC_3_743, output_MAC_3_744, output_MAC_3_745, output_MAC_3_746, output_MAC_3_747, output_MAC_3_748, output_MAC_3_749, 
		output_MAC_3_750, output_MAC_3_751, output_MAC_3_752, output_MAC_3_753, output_MAC_3_754, output_MAC_3_755, output_MAC_3_756, output_MAC_3_757, output_MAC_3_758, output_MAC_3_759, 
		output_MAC_3_760, output_MAC_3_761, output_MAC_3_762, output_MAC_3_763, output_MAC_3_764, output_MAC_3_765, output_MAC_3_766, output_MAC_3_767: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_4_0, output_MAC_4_1, output_MAC_4_2, output_MAC_4_3, output_MAC_4_4, output_MAC_4_5, output_MAC_4_6, output_MAC_4_7, output_MAC_4_8, output_MAC_4_9, 
		output_MAC_4_10, output_MAC_4_11, output_MAC_4_12, output_MAC_4_13, output_MAC_4_14, output_MAC_4_15, output_MAC_4_16, output_MAC_4_17, output_MAC_4_18, output_MAC_4_19, 
		output_MAC_4_20, output_MAC_4_21, output_MAC_4_22, output_MAC_4_23, output_MAC_4_24, output_MAC_4_25, output_MAC_4_26, output_MAC_4_27, output_MAC_4_28, output_MAC_4_29, 
		output_MAC_4_30, output_MAC_4_31, output_MAC_4_32, output_MAC_4_33, output_MAC_4_34, output_MAC_4_35, output_MAC_4_36, output_MAC_4_37, output_MAC_4_38, output_MAC_4_39, 
		output_MAC_4_40, output_MAC_4_41, output_MAC_4_42, output_MAC_4_43, output_MAC_4_44, output_MAC_4_45, output_MAC_4_46, output_MAC_4_47, output_MAC_4_48, output_MAC_4_49, 
		output_MAC_4_50, output_MAC_4_51, output_MAC_4_52, output_MAC_4_53, output_MAC_4_54, output_MAC_4_55, output_MAC_4_56, output_MAC_4_57, output_MAC_4_58, output_MAC_4_59, 
		output_MAC_4_60, output_MAC_4_61, output_MAC_4_62, output_MAC_4_63, output_MAC_4_64, output_MAC_4_65, output_MAC_4_66, output_MAC_4_67, output_MAC_4_68, output_MAC_4_69, 
		output_MAC_4_70, output_MAC_4_71, output_MAC_4_72, output_MAC_4_73, output_MAC_4_74, output_MAC_4_75, output_MAC_4_76, output_MAC_4_77, output_MAC_4_78, output_MAC_4_79, 
		output_MAC_4_80, output_MAC_4_81, output_MAC_4_82, output_MAC_4_83, output_MAC_4_84, output_MAC_4_85, output_MAC_4_86, output_MAC_4_87, output_MAC_4_88, output_MAC_4_89, 
		output_MAC_4_90, output_MAC_4_91, output_MAC_4_92, output_MAC_4_93, output_MAC_4_94, output_MAC_4_95, output_MAC_4_96, output_MAC_4_97, output_MAC_4_98, output_MAC_4_99, 
		output_MAC_4_100, output_MAC_4_101, output_MAC_4_102, output_MAC_4_103, output_MAC_4_104, output_MAC_4_105, output_MAC_4_106, output_MAC_4_107, output_MAC_4_108, output_MAC_4_109, 
		output_MAC_4_110, output_MAC_4_111, output_MAC_4_112, output_MAC_4_113, output_MAC_4_114, output_MAC_4_115, output_MAC_4_116, output_MAC_4_117, output_MAC_4_118, output_MAC_4_119, 
		output_MAC_4_120, output_MAC_4_121, output_MAC_4_122, output_MAC_4_123, output_MAC_4_124, output_MAC_4_125, output_MAC_4_126, output_MAC_4_127, output_MAC_4_128, output_MAC_4_129, 
		output_MAC_4_130, output_MAC_4_131, output_MAC_4_132, output_MAC_4_133, output_MAC_4_134, output_MAC_4_135, output_MAC_4_136, output_MAC_4_137, output_MAC_4_138, output_MAC_4_139, 
		output_MAC_4_140, output_MAC_4_141, output_MAC_4_142, output_MAC_4_143, output_MAC_4_144, output_MAC_4_145, output_MAC_4_146, output_MAC_4_147, output_MAC_4_148, output_MAC_4_149, 
		output_MAC_4_150, output_MAC_4_151, output_MAC_4_152, output_MAC_4_153, output_MAC_4_154, output_MAC_4_155, output_MAC_4_156, output_MAC_4_157, output_MAC_4_158, output_MAC_4_159, 
		output_MAC_4_160, output_MAC_4_161, output_MAC_4_162, output_MAC_4_163, output_MAC_4_164, output_MAC_4_165, output_MAC_4_166, output_MAC_4_167, output_MAC_4_168, output_MAC_4_169, 
		output_MAC_4_170, output_MAC_4_171, output_MAC_4_172, output_MAC_4_173, output_MAC_4_174, output_MAC_4_175, output_MAC_4_176, output_MAC_4_177, output_MAC_4_178, output_MAC_4_179, 
		output_MAC_4_180, output_MAC_4_181, output_MAC_4_182, output_MAC_4_183, output_MAC_4_184, output_MAC_4_185, output_MAC_4_186, output_MAC_4_187, output_MAC_4_188, output_MAC_4_189, 
		output_MAC_4_190, output_MAC_4_191, output_MAC_4_192, output_MAC_4_193, output_MAC_4_194, output_MAC_4_195, output_MAC_4_196, output_MAC_4_197, output_MAC_4_198, output_MAC_4_199, 
		output_MAC_4_200, output_MAC_4_201, output_MAC_4_202, output_MAC_4_203, output_MAC_4_204, output_MAC_4_205, output_MAC_4_206, output_MAC_4_207, output_MAC_4_208, output_MAC_4_209, 
		output_MAC_4_210, output_MAC_4_211, output_MAC_4_212, output_MAC_4_213, output_MAC_4_214, output_MAC_4_215, output_MAC_4_216, output_MAC_4_217, output_MAC_4_218, output_MAC_4_219, 
		output_MAC_4_220, output_MAC_4_221, output_MAC_4_222, output_MAC_4_223, output_MAC_4_224, output_MAC_4_225, output_MAC_4_226, output_MAC_4_227, output_MAC_4_228, output_MAC_4_229, 
		output_MAC_4_230, output_MAC_4_231, output_MAC_4_232, output_MAC_4_233, output_MAC_4_234, output_MAC_4_235, output_MAC_4_236, output_MAC_4_237, output_MAC_4_238, output_MAC_4_239, 
		output_MAC_4_240, output_MAC_4_241, output_MAC_4_242, output_MAC_4_243, output_MAC_4_244, output_MAC_4_245, output_MAC_4_246, output_MAC_4_247, output_MAC_4_248, output_MAC_4_249, 
		output_MAC_4_250, output_MAC_4_251, output_MAC_4_252, output_MAC_4_253, output_MAC_4_254, output_MAC_4_255, output_MAC_4_256, output_MAC_4_257, output_MAC_4_258, output_MAC_4_259, 
		output_MAC_4_260, output_MAC_4_261, output_MAC_4_262, output_MAC_4_263, output_MAC_4_264, output_MAC_4_265, output_MAC_4_266, output_MAC_4_267, output_MAC_4_268, output_MAC_4_269, 
		output_MAC_4_270, output_MAC_4_271, output_MAC_4_272, output_MAC_4_273, output_MAC_4_274, output_MAC_4_275, output_MAC_4_276, output_MAC_4_277, output_MAC_4_278, output_MAC_4_279, 
		output_MAC_4_280, output_MAC_4_281, output_MAC_4_282, output_MAC_4_283, output_MAC_4_284, output_MAC_4_285, output_MAC_4_286, output_MAC_4_287, output_MAC_4_288, output_MAC_4_289, 
		output_MAC_4_290, output_MAC_4_291, output_MAC_4_292, output_MAC_4_293, output_MAC_4_294, output_MAC_4_295, output_MAC_4_296, output_MAC_4_297, output_MAC_4_298, output_MAC_4_299, 
		output_MAC_4_300, output_MAC_4_301, output_MAC_4_302, output_MAC_4_303, output_MAC_4_304, output_MAC_4_305, output_MAC_4_306, output_MAC_4_307, output_MAC_4_308, output_MAC_4_309, 
		output_MAC_4_310, output_MAC_4_311, output_MAC_4_312, output_MAC_4_313, output_MAC_4_314, output_MAC_4_315, output_MAC_4_316, output_MAC_4_317, output_MAC_4_318, output_MAC_4_319, 
		output_MAC_4_320, output_MAC_4_321, output_MAC_4_322, output_MAC_4_323, output_MAC_4_324, output_MAC_4_325, output_MAC_4_326, output_MAC_4_327, output_MAC_4_328, output_MAC_4_329, 
		output_MAC_4_330, output_MAC_4_331, output_MAC_4_332, output_MAC_4_333, output_MAC_4_334, output_MAC_4_335, output_MAC_4_336, output_MAC_4_337, output_MAC_4_338, output_MAC_4_339, 
		output_MAC_4_340, output_MAC_4_341, output_MAC_4_342, output_MAC_4_343, output_MAC_4_344, output_MAC_4_345, output_MAC_4_346, output_MAC_4_347, output_MAC_4_348, output_MAC_4_349, 
		output_MAC_4_350, output_MAC_4_351, output_MAC_4_352, output_MAC_4_353, output_MAC_4_354, output_MAC_4_355, output_MAC_4_356, output_MAC_4_357, output_MAC_4_358, output_MAC_4_359, 
		output_MAC_4_360, output_MAC_4_361, output_MAC_4_362, output_MAC_4_363, output_MAC_4_364, output_MAC_4_365, output_MAC_4_366, output_MAC_4_367, output_MAC_4_368, output_MAC_4_369, 
		output_MAC_4_370, output_MAC_4_371, output_MAC_4_372, output_MAC_4_373, output_MAC_4_374, output_MAC_4_375, output_MAC_4_376, output_MAC_4_377, output_MAC_4_378, output_MAC_4_379, 
		output_MAC_4_380, output_MAC_4_381, output_MAC_4_382, output_MAC_4_383, output_MAC_4_384, output_MAC_4_385, output_MAC_4_386, output_MAC_4_387, output_MAC_4_388, output_MAC_4_389, 
		output_MAC_4_390, output_MAC_4_391, output_MAC_4_392, output_MAC_4_393, output_MAC_4_394, output_MAC_4_395, output_MAC_4_396, output_MAC_4_397, output_MAC_4_398, output_MAC_4_399, 
		output_MAC_4_400, output_MAC_4_401, output_MAC_4_402, output_MAC_4_403, output_MAC_4_404, output_MAC_4_405, output_MAC_4_406, output_MAC_4_407, output_MAC_4_408, output_MAC_4_409, 
		output_MAC_4_410, output_MAC_4_411, output_MAC_4_412, output_MAC_4_413, output_MAC_4_414, output_MAC_4_415, output_MAC_4_416, output_MAC_4_417, output_MAC_4_418, output_MAC_4_419, 
		output_MAC_4_420, output_MAC_4_421, output_MAC_4_422, output_MAC_4_423, output_MAC_4_424, output_MAC_4_425, output_MAC_4_426, output_MAC_4_427, output_MAC_4_428, output_MAC_4_429, 
		output_MAC_4_430, output_MAC_4_431, output_MAC_4_432, output_MAC_4_433, output_MAC_4_434, output_MAC_4_435, output_MAC_4_436, output_MAC_4_437, output_MAC_4_438, output_MAC_4_439, 
		output_MAC_4_440, output_MAC_4_441, output_MAC_4_442, output_MAC_4_443, output_MAC_4_444, output_MAC_4_445, output_MAC_4_446, output_MAC_4_447, output_MAC_4_448, output_MAC_4_449, 
		output_MAC_4_450, output_MAC_4_451, output_MAC_4_452, output_MAC_4_453, output_MAC_4_454, output_MAC_4_455, output_MAC_4_456, output_MAC_4_457, output_MAC_4_458, output_MAC_4_459, 
		output_MAC_4_460, output_MAC_4_461, output_MAC_4_462, output_MAC_4_463, output_MAC_4_464, output_MAC_4_465, output_MAC_4_466, output_MAC_4_467, output_MAC_4_468, output_MAC_4_469, 
		output_MAC_4_470, output_MAC_4_471, output_MAC_4_472, output_MAC_4_473, output_MAC_4_474, output_MAC_4_475, output_MAC_4_476, output_MAC_4_477, output_MAC_4_478, output_MAC_4_479, 
		output_MAC_4_480, output_MAC_4_481, output_MAC_4_482, output_MAC_4_483, output_MAC_4_484, output_MAC_4_485, output_MAC_4_486, output_MAC_4_487, output_MAC_4_488, output_MAC_4_489, 
		output_MAC_4_490, output_MAC_4_491, output_MAC_4_492, output_MAC_4_493, output_MAC_4_494, output_MAC_4_495, output_MAC_4_496, output_MAC_4_497, output_MAC_4_498, output_MAC_4_499, 
		output_MAC_4_500, output_MAC_4_501, output_MAC_4_502, output_MAC_4_503, output_MAC_4_504, output_MAC_4_505, output_MAC_4_506, output_MAC_4_507, output_MAC_4_508, output_MAC_4_509, 
		output_MAC_4_510, output_MAC_4_511, output_MAC_4_512, output_MAC_4_513, output_MAC_4_514, output_MAC_4_515, output_MAC_4_516, output_MAC_4_517, output_MAC_4_518, output_MAC_4_519, 
		output_MAC_4_520, output_MAC_4_521, output_MAC_4_522, output_MAC_4_523, output_MAC_4_524, output_MAC_4_525, output_MAC_4_526, output_MAC_4_527, output_MAC_4_528, output_MAC_4_529, 
		output_MAC_4_530, output_MAC_4_531, output_MAC_4_532, output_MAC_4_533, output_MAC_4_534, output_MAC_4_535, output_MAC_4_536, output_MAC_4_537, output_MAC_4_538, output_MAC_4_539, 
		output_MAC_4_540, output_MAC_4_541, output_MAC_4_542, output_MAC_4_543, output_MAC_4_544, output_MAC_4_545, output_MAC_4_546, output_MAC_4_547, output_MAC_4_548, output_MAC_4_549, 
		output_MAC_4_550, output_MAC_4_551, output_MAC_4_552, output_MAC_4_553, output_MAC_4_554, output_MAC_4_555, output_MAC_4_556, output_MAC_4_557, output_MAC_4_558, output_MAC_4_559, 
		output_MAC_4_560, output_MAC_4_561, output_MAC_4_562, output_MAC_4_563, output_MAC_4_564, output_MAC_4_565, output_MAC_4_566, output_MAC_4_567, output_MAC_4_568, output_MAC_4_569, 
		output_MAC_4_570, output_MAC_4_571, output_MAC_4_572, output_MAC_4_573, output_MAC_4_574, output_MAC_4_575, output_MAC_4_576, output_MAC_4_577, output_MAC_4_578, output_MAC_4_579, 
		output_MAC_4_580, output_MAC_4_581, output_MAC_4_582, output_MAC_4_583, output_MAC_4_584, output_MAC_4_585, output_MAC_4_586, output_MAC_4_587, output_MAC_4_588, output_MAC_4_589, 
		output_MAC_4_590, output_MAC_4_591, output_MAC_4_592, output_MAC_4_593, output_MAC_4_594, output_MAC_4_595, output_MAC_4_596, output_MAC_4_597, output_MAC_4_598, output_MAC_4_599, 
		output_MAC_4_600, output_MAC_4_601, output_MAC_4_602, output_MAC_4_603, output_MAC_4_604, output_MAC_4_605, output_MAC_4_606, output_MAC_4_607, output_MAC_4_608, output_MAC_4_609, 
		output_MAC_4_610, output_MAC_4_611, output_MAC_4_612, output_MAC_4_613, output_MAC_4_614, output_MAC_4_615, output_MAC_4_616, output_MAC_4_617, output_MAC_4_618, output_MAC_4_619, 
		output_MAC_4_620, output_MAC_4_621, output_MAC_4_622, output_MAC_4_623, output_MAC_4_624, output_MAC_4_625, output_MAC_4_626, output_MAC_4_627, output_MAC_4_628, output_MAC_4_629, 
		output_MAC_4_630, output_MAC_4_631, output_MAC_4_632, output_MAC_4_633, output_MAC_4_634, output_MAC_4_635, output_MAC_4_636, output_MAC_4_637, output_MAC_4_638, output_MAC_4_639, 
		output_MAC_4_640, output_MAC_4_641, output_MAC_4_642, output_MAC_4_643, output_MAC_4_644, output_MAC_4_645, output_MAC_4_646, output_MAC_4_647, output_MAC_4_648, output_MAC_4_649, 
		output_MAC_4_650, output_MAC_4_651, output_MAC_4_652, output_MAC_4_653, output_MAC_4_654, output_MAC_4_655, output_MAC_4_656, output_MAC_4_657, output_MAC_4_658, output_MAC_4_659, 
		output_MAC_4_660, output_MAC_4_661, output_MAC_4_662, output_MAC_4_663, output_MAC_4_664, output_MAC_4_665, output_MAC_4_666, output_MAC_4_667, output_MAC_4_668, output_MAC_4_669, 
		output_MAC_4_670, output_MAC_4_671, output_MAC_4_672, output_MAC_4_673, output_MAC_4_674, output_MAC_4_675, output_MAC_4_676, output_MAC_4_677, output_MAC_4_678, output_MAC_4_679, 
		output_MAC_4_680, output_MAC_4_681, output_MAC_4_682, output_MAC_4_683, output_MAC_4_684, output_MAC_4_685, output_MAC_4_686, output_MAC_4_687, output_MAC_4_688, output_MAC_4_689, 
		output_MAC_4_690, output_MAC_4_691, output_MAC_4_692, output_MAC_4_693, output_MAC_4_694, output_MAC_4_695, output_MAC_4_696, output_MAC_4_697, output_MAC_4_698, output_MAC_4_699, 
		output_MAC_4_700, output_MAC_4_701, output_MAC_4_702, output_MAC_4_703, output_MAC_4_704, output_MAC_4_705, output_MAC_4_706, output_MAC_4_707, output_MAC_4_708, output_MAC_4_709, 
		output_MAC_4_710, output_MAC_4_711, output_MAC_4_712, output_MAC_4_713, output_MAC_4_714, output_MAC_4_715, output_MAC_4_716, output_MAC_4_717, output_MAC_4_718, output_MAC_4_719, 
		output_MAC_4_720, output_MAC_4_721, output_MAC_4_722, output_MAC_4_723, output_MAC_4_724, output_MAC_4_725, output_MAC_4_726, output_MAC_4_727, output_MAC_4_728, output_MAC_4_729, 
		output_MAC_4_730, output_MAC_4_731, output_MAC_4_732, output_MAC_4_733, output_MAC_4_734, output_MAC_4_735, output_MAC_4_736, output_MAC_4_737, output_MAC_4_738, output_MAC_4_739, 
		output_MAC_4_740, output_MAC_4_741, output_MAC_4_742, output_MAC_4_743, output_MAC_4_744, output_MAC_4_745, output_MAC_4_746, output_MAC_4_747, output_MAC_4_748, output_MAC_4_749, 
		output_MAC_4_750, output_MAC_4_751, output_MAC_4_752, output_MAC_4_753, output_MAC_4_754, output_MAC_4_755, output_MAC_4_756, output_MAC_4_757, output_MAC_4_758, output_MAC_4_759, 
		output_MAC_4_760, output_MAC_4_761, output_MAC_4_762, output_MAC_4_763, output_MAC_4_764, output_MAC_4_765, output_MAC_4_766, output_MAC_4_767: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_5_0, output_MAC_5_1, output_MAC_5_2, output_MAC_5_3, output_MAC_5_4, output_MAC_5_5, output_MAC_5_6, output_MAC_5_7, output_MAC_5_8, output_MAC_5_9, 
		output_MAC_5_10, output_MAC_5_11, output_MAC_5_12, output_MAC_5_13, output_MAC_5_14, output_MAC_5_15, output_MAC_5_16, output_MAC_5_17, output_MAC_5_18, output_MAC_5_19, 
		output_MAC_5_20, output_MAC_5_21, output_MAC_5_22, output_MAC_5_23, output_MAC_5_24, output_MAC_5_25, output_MAC_5_26, output_MAC_5_27, output_MAC_5_28, output_MAC_5_29, 
		output_MAC_5_30, output_MAC_5_31, output_MAC_5_32, output_MAC_5_33, output_MAC_5_34, output_MAC_5_35, output_MAC_5_36, output_MAC_5_37, output_MAC_5_38, output_MAC_5_39, 
		output_MAC_5_40, output_MAC_5_41, output_MAC_5_42, output_MAC_5_43, output_MAC_5_44, output_MAC_5_45, output_MAC_5_46, output_MAC_5_47, output_MAC_5_48, output_MAC_5_49, 
		output_MAC_5_50, output_MAC_5_51, output_MAC_5_52, output_MAC_5_53, output_MAC_5_54, output_MAC_5_55, output_MAC_5_56, output_MAC_5_57, output_MAC_5_58, output_MAC_5_59, 
		output_MAC_5_60, output_MAC_5_61, output_MAC_5_62, output_MAC_5_63, output_MAC_5_64, output_MAC_5_65, output_MAC_5_66, output_MAC_5_67, output_MAC_5_68, output_MAC_5_69, 
		output_MAC_5_70, output_MAC_5_71, output_MAC_5_72, output_MAC_5_73, output_MAC_5_74, output_MAC_5_75, output_MAC_5_76, output_MAC_5_77, output_MAC_5_78, output_MAC_5_79, 
		output_MAC_5_80, output_MAC_5_81, output_MAC_5_82, output_MAC_5_83, output_MAC_5_84, output_MAC_5_85, output_MAC_5_86, output_MAC_5_87, output_MAC_5_88, output_MAC_5_89, 
		output_MAC_5_90, output_MAC_5_91, output_MAC_5_92, output_MAC_5_93, output_MAC_5_94, output_MAC_5_95, output_MAC_5_96, output_MAC_5_97, output_MAC_5_98, output_MAC_5_99, 
		output_MAC_5_100, output_MAC_5_101, output_MAC_5_102, output_MAC_5_103, output_MAC_5_104, output_MAC_5_105, output_MAC_5_106, output_MAC_5_107, output_MAC_5_108, output_MAC_5_109, 
		output_MAC_5_110, output_MAC_5_111, output_MAC_5_112, output_MAC_5_113, output_MAC_5_114, output_MAC_5_115, output_MAC_5_116, output_MAC_5_117, output_MAC_5_118, output_MAC_5_119, 
		output_MAC_5_120, output_MAC_5_121, output_MAC_5_122, output_MAC_5_123, output_MAC_5_124, output_MAC_5_125, output_MAC_5_126, output_MAC_5_127, output_MAC_5_128, output_MAC_5_129, 
		output_MAC_5_130, output_MAC_5_131, output_MAC_5_132, output_MAC_5_133, output_MAC_5_134, output_MAC_5_135, output_MAC_5_136, output_MAC_5_137, output_MAC_5_138, output_MAC_5_139, 
		output_MAC_5_140, output_MAC_5_141, output_MAC_5_142, output_MAC_5_143, output_MAC_5_144, output_MAC_5_145, output_MAC_5_146, output_MAC_5_147, output_MAC_5_148, output_MAC_5_149, 
		output_MAC_5_150, output_MAC_5_151, output_MAC_5_152, output_MAC_5_153, output_MAC_5_154, output_MAC_5_155, output_MAC_5_156, output_MAC_5_157, output_MAC_5_158, output_MAC_5_159, 
		output_MAC_5_160, output_MAC_5_161, output_MAC_5_162, output_MAC_5_163, output_MAC_5_164, output_MAC_5_165, output_MAC_5_166, output_MAC_5_167, output_MAC_5_168, output_MAC_5_169, 
		output_MAC_5_170, output_MAC_5_171, output_MAC_5_172, output_MAC_5_173, output_MAC_5_174, output_MAC_5_175, output_MAC_5_176, output_MAC_5_177, output_MAC_5_178, output_MAC_5_179, 
		output_MAC_5_180, output_MAC_5_181, output_MAC_5_182, output_MAC_5_183, output_MAC_5_184, output_MAC_5_185, output_MAC_5_186, output_MAC_5_187, output_MAC_5_188, output_MAC_5_189, 
		output_MAC_5_190, output_MAC_5_191, output_MAC_5_192, output_MAC_5_193, output_MAC_5_194, output_MAC_5_195, output_MAC_5_196, output_MAC_5_197, output_MAC_5_198, output_MAC_5_199, 
		output_MAC_5_200, output_MAC_5_201, output_MAC_5_202, output_MAC_5_203, output_MAC_5_204, output_MAC_5_205, output_MAC_5_206, output_MAC_5_207, output_MAC_5_208, output_MAC_5_209, 
		output_MAC_5_210, output_MAC_5_211, output_MAC_5_212, output_MAC_5_213, output_MAC_5_214, output_MAC_5_215, output_MAC_5_216, output_MAC_5_217, output_MAC_5_218, output_MAC_5_219, 
		output_MAC_5_220, output_MAC_5_221, output_MAC_5_222, output_MAC_5_223, output_MAC_5_224, output_MAC_5_225, output_MAC_5_226, output_MAC_5_227, output_MAC_5_228, output_MAC_5_229, 
		output_MAC_5_230, output_MAC_5_231, output_MAC_5_232, output_MAC_5_233, output_MAC_5_234, output_MAC_5_235, output_MAC_5_236, output_MAC_5_237, output_MAC_5_238, output_MAC_5_239, 
		output_MAC_5_240, output_MAC_5_241, output_MAC_5_242, output_MAC_5_243, output_MAC_5_244, output_MAC_5_245, output_MAC_5_246, output_MAC_5_247, output_MAC_5_248, output_MAC_5_249, 
		output_MAC_5_250, output_MAC_5_251, output_MAC_5_252, output_MAC_5_253, output_MAC_5_254, output_MAC_5_255, output_MAC_5_256, output_MAC_5_257, output_MAC_5_258, output_MAC_5_259, 
		output_MAC_5_260, output_MAC_5_261, output_MAC_5_262, output_MAC_5_263, output_MAC_5_264, output_MAC_5_265, output_MAC_5_266, output_MAC_5_267, output_MAC_5_268, output_MAC_5_269, 
		output_MAC_5_270, output_MAC_5_271, output_MAC_5_272, output_MAC_5_273, output_MAC_5_274, output_MAC_5_275, output_MAC_5_276, output_MAC_5_277, output_MAC_5_278, output_MAC_5_279, 
		output_MAC_5_280, output_MAC_5_281, output_MAC_5_282, output_MAC_5_283, output_MAC_5_284, output_MAC_5_285, output_MAC_5_286, output_MAC_5_287, output_MAC_5_288, output_MAC_5_289, 
		output_MAC_5_290, output_MAC_5_291, output_MAC_5_292, output_MAC_5_293, output_MAC_5_294, output_MAC_5_295, output_MAC_5_296, output_MAC_5_297, output_MAC_5_298, output_MAC_5_299, 
		output_MAC_5_300, output_MAC_5_301, output_MAC_5_302, output_MAC_5_303, output_MAC_5_304, output_MAC_5_305, output_MAC_5_306, output_MAC_5_307, output_MAC_5_308, output_MAC_5_309, 
		output_MAC_5_310, output_MAC_5_311, output_MAC_5_312, output_MAC_5_313, output_MAC_5_314, output_MAC_5_315, output_MAC_5_316, output_MAC_5_317, output_MAC_5_318, output_MAC_5_319, 
		output_MAC_5_320, output_MAC_5_321, output_MAC_5_322, output_MAC_5_323, output_MAC_5_324, output_MAC_5_325, output_MAC_5_326, output_MAC_5_327, output_MAC_5_328, output_MAC_5_329, 
		output_MAC_5_330, output_MAC_5_331, output_MAC_5_332, output_MAC_5_333, output_MAC_5_334, output_MAC_5_335, output_MAC_5_336, output_MAC_5_337, output_MAC_5_338, output_MAC_5_339, 
		output_MAC_5_340, output_MAC_5_341, output_MAC_5_342, output_MAC_5_343, output_MAC_5_344, output_MAC_5_345, output_MAC_5_346, output_MAC_5_347, output_MAC_5_348, output_MAC_5_349, 
		output_MAC_5_350, output_MAC_5_351, output_MAC_5_352, output_MAC_5_353, output_MAC_5_354, output_MAC_5_355, output_MAC_5_356, output_MAC_5_357, output_MAC_5_358, output_MAC_5_359, 
		output_MAC_5_360, output_MAC_5_361, output_MAC_5_362, output_MAC_5_363, output_MAC_5_364, output_MAC_5_365, output_MAC_5_366, output_MAC_5_367, output_MAC_5_368, output_MAC_5_369, 
		output_MAC_5_370, output_MAC_5_371, output_MAC_5_372, output_MAC_5_373, output_MAC_5_374, output_MAC_5_375, output_MAC_5_376, output_MAC_5_377, output_MAC_5_378, output_MAC_5_379, 
		output_MAC_5_380, output_MAC_5_381, output_MAC_5_382, output_MAC_5_383, output_MAC_5_384, output_MAC_5_385, output_MAC_5_386, output_MAC_5_387, output_MAC_5_388, output_MAC_5_389, 
		output_MAC_5_390, output_MAC_5_391, output_MAC_5_392, output_MAC_5_393, output_MAC_5_394, output_MAC_5_395, output_MAC_5_396, output_MAC_5_397, output_MAC_5_398, output_MAC_5_399, 
		output_MAC_5_400, output_MAC_5_401, output_MAC_5_402, output_MAC_5_403, output_MAC_5_404, output_MAC_5_405, output_MAC_5_406, output_MAC_5_407, output_MAC_5_408, output_MAC_5_409, 
		output_MAC_5_410, output_MAC_5_411, output_MAC_5_412, output_MAC_5_413, output_MAC_5_414, output_MAC_5_415, output_MAC_5_416, output_MAC_5_417, output_MAC_5_418, output_MAC_5_419, 
		output_MAC_5_420, output_MAC_5_421, output_MAC_5_422, output_MAC_5_423, output_MAC_5_424, output_MAC_5_425, output_MAC_5_426, output_MAC_5_427, output_MAC_5_428, output_MAC_5_429, 
		output_MAC_5_430, output_MAC_5_431, output_MAC_5_432, output_MAC_5_433, output_MAC_5_434, output_MAC_5_435, output_MAC_5_436, output_MAC_5_437, output_MAC_5_438, output_MAC_5_439, 
		output_MAC_5_440, output_MAC_5_441, output_MAC_5_442, output_MAC_5_443, output_MAC_5_444, output_MAC_5_445, output_MAC_5_446, output_MAC_5_447, output_MAC_5_448, output_MAC_5_449, 
		output_MAC_5_450, output_MAC_5_451, output_MAC_5_452, output_MAC_5_453, output_MAC_5_454, output_MAC_5_455, output_MAC_5_456, output_MAC_5_457, output_MAC_5_458, output_MAC_5_459, 
		output_MAC_5_460, output_MAC_5_461, output_MAC_5_462, output_MAC_5_463, output_MAC_5_464, output_MAC_5_465, output_MAC_5_466, output_MAC_5_467, output_MAC_5_468, output_MAC_5_469, 
		output_MAC_5_470, output_MAC_5_471, output_MAC_5_472, output_MAC_5_473, output_MAC_5_474, output_MAC_5_475, output_MAC_5_476, output_MAC_5_477, output_MAC_5_478, output_MAC_5_479, 
		output_MAC_5_480, output_MAC_5_481, output_MAC_5_482, output_MAC_5_483, output_MAC_5_484, output_MAC_5_485, output_MAC_5_486, output_MAC_5_487, output_MAC_5_488, output_MAC_5_489, 
		output_MAC_5_490, output_MAC_5_491, output_MAC_5_492, output_MAC_5_493, output_MAC_5_494, output_MAC_5_495, output_MAC_5_496, output_MAC_5_497, output_MAC_5_498, output_MAC_5_499, 
		output_MAC_5_500, output_MAC_5_501, output_MAC_5_502, output_MAC_5_503, output_MAC_5_504, output_MAC_5_505, output_MAC_5_506, output_MAC_5_507, output_MAC_5_508, output_MAC_5_509, 
		output_MAC_5_510, output_MAC_5_511, output_MAC_5_512, output_MAC_5_513, output_MAC_5_514, output_MAC_5_515, output_MAC_5_516, output_MAC_5_517, output_MAC_5_518, output_MAC_5_519, 
		output_MAC_5_520, output_MAC_5_521, output_MAC_5_522, output_MAC_5_523, output_MAC_5_524, output_MAC_5_525, output_MAC_5_526, output_MAC_5_527, output_MAC_5_528, output_MAC_5_529, 
		output_MAC_5_530, output_MAC_5_531, output_MAC_5_532, output_MAC_5_533, output_MAC_5_534, output_MAC_5_535, output_MAC_5_536, output_MAC_5_537, output_MAC_5_538, output_MAC_5_539, 
		output_MAC_5_540, output_MAC_5_541, output_MAC_5_542, output_MAC_5_543, output_MAC_5_544, output_MAC_5_545, output_MAC_5_546, output_MAC_5_547, output_MAC_5_548, output_MAC_5_549, 
		output_MAC_5_550, output_MAC_5_551, output_MAC_5_552, output_MAC_5_553, output_MAC_5_554, output_MAC_5_555, output_MAC_5_556, output_MAC_5_557, output_MAC_5_558, output_MAC_5_559, 
		output_MAC_5_560, output_MAC_5_561, output_MAC_5_562, output_MAC_5_563, output_MAC_5_564, output_MAC_5_565, output_MAC_5_566, output_MAC_5_567, output_MAC_5_568, output_MAC_5_569, 
		output_MAC_5_570, output_MAC_5_571, output_MAC_5_572, output_MAC_5_573, output_MAC_5_574, output_MAC_5_575, output_MAC_5_576, output_MAC_5_577, output_MAC_5_578, output_MAC_5_579, 
		output_MAC_5_580, output_MAC_5_581, output_MAC_5_582, output_MAC_5_583, output_MAC_5_584, output_MAC_5_585, output_MAC_5_586, output_MAC_5_587, output_MAC_5_588, output_MAC_5_589, 
		output_MAC_5_590, output_MAC_5_591, output_MAC_5_592, output_MAC_5_593, output_MAC_5_594, output_MAC_5_595, output_MAC_5_596, output_MAC_5_597, output_MAC_5_598, output_MAC_5_599, 
		output_MAC_5_600, output_MAC_5_601, output_MAC_5_602, output_MAC_5_603, output_MAC_5_604, output_MAC_5_605, output_MAC_5_606, output_MAC_5_607, output_MAC_5_608, output_MAC_5_609, 
		output_MAC_5_610, output_MAC_5_611, output_MAC_5_612, output_MAC_5_613, output_MAC_5_614, output_MAC_5_615, output_MAC_5_616, output_MAC_5_617, output_MAC_5_618, output_MAC_5_619, 
		output_MAC_5_620, output_MAC_5_621, output_MAC_5_622, output_MAC_5_623, output_MAC_5_624, output_MAC_5_625, output_MAC_5_626, output_MAC_5_627, output_MAC_5_628, output_MAC_5_629, 
		output_MAC_5_630, output_MAC_5_631, output_MAC_5_632, output_MAC_5_633, output_MAC_5_634, output_MAC_5_635, output_MAC_5_636, output_MAC_5_637, output_MAC_5_638, output_MAC_5_639, 
		output_MAC_5_640, output_MAC_5_641, output_MAC_5_642, output_MAC_5_643, output_MAC_5_644, output_MAC_5_645, output_MAC_5_646, output_MAC_5_647, output_MAC_5_648, output_MAC_5_649, 
		output_MAC_5_650, output_MAC_5_651, output_MAC_5_652, output_MAC_5_653, output_MAC_5_654, output_MAC_5_655, output_MAC_5_656, output_MAC_5_657, output_MAC_5_658, output_MAC_5_659, 
		output_MAC_5_660, output_MAC_5_661, output_MAC_5_662, output_MAC_5_663, output_MAC_5_664, output_MAC_5_665, output_MAC_5_666, output_MAC_5_667, output_MAC_5_668, output_MAC_5_669, 
		output_MAC_5_670, output_MAC_5_671, output_MAC_5_672, output_MAC_5_673, output_MAC_5_674, output_MAC_5_675, output_MAC_5_676, output_MAC_5_677, output_MAC_5_678, output_MAC_5_679, 
		output_MAC_5_680, output_MAC_5_681, output_MAC_5_682, output_MAC_5_683, output_MAC_5_684, output_MAC_5_685, output_MAC_5_686, output_MAC_5_687, output_MAC_5_688, output_MAC_5_689, 
		output_MAC_5_690, output_MAC_5_691, output_MAC_5_692, output_MAC_5_693, output_MAC_5_694, output_MAC_5_695, output_MAC_5_696, output_MAC_5_697, output_MAC_5_698, output_MAC_5_699, 
		output_MAC_5_700, output_MAC_5_701, output_MAC_5_702, output_MAC_5_703, output_MAC_5_704, output_MAC_5_705, output_MAC_5_706, output_MAC_5_707, output_MAC_5_708, output_MAC_5_709, 
		output_MAC_5_710, output_MAC_5_711, output_MAC_5_712, output_MAC_5_713, output_MAC_5_714, output_MAC_5_715, output_MAC_5_716, output_MAC_5_717, output_MAC_5_718, output_MAC_5_719, 
		output_MAC_5_720, output_MAC_5_721, output_MAC_5_722, output_MAC_5_723, output_MAC_5_724, output_MAC_5_725, output_MAC_5_726, output_MAC_5_727, output_MAC_5_728, output_MAC_5_729, 
		output_MAC_5_730, output_MAC_5_731, output_MAC_5_732, output_MAC_5_733, output_MAC_5_734, output_MAC_5_735, output_MAC_5_736, output_MAC_5_737, output_MAC_5_738, output_MAC_5_739, 
		output_MAC_5_740, output_MAC_5_741, output_MAC_5_742, output_MAC_5_743, output_MAC_5_744, output_MAC_5_745, output_MAC_5_746, output_MAC_5_747, output_MAC_5_748, output_MAC_5_749, 
		output_MAC_5_750, output_MAC_5_751, output_MAC_5_752, output_MAC_5_753, output_MAC_5_754, output_MAC_5_755, output_MAC_5_756, output_MAC_5_757, output_MAC_5_758, output_MAC_5_759, 
		output_MAC_5_760, output_MAC_5_761, output_MAC_5_762, output_MAC_5_763, output_MAC_5_764, output_MAC_5_765, output_MAC_5_766, output_MAC_5_767: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_6_0, output_MAC_6_1, output_MAC_6_2, output_MAC_6_3, output_MAC_6_4, output_MAC_6_5, output_MAC_6_6, output_MAC_6_7, output_MAC_6_8, output_MAC_6_9, 
		output_MAC_6_10, output_MAC_6_11, output_MAC_6_12, output_MAC_6_13, output_MAC_6_14, output_MAC_6_15, output_MAC_6_16, output_MAC_6_17, output_MAC_6_18, output_MAC_6_19, 
		output_MAC_6_20, output_MAC_6_21, output_MAC_6_22, output_MAC_6_23, output_MAC_6_24, output_MAC_6_25, output_MAC_6_26, output_MAC_6_27, output_MAC_6_28, output_MAC_6_29, 
		output_MAC_6_30, output_MAC_6_31, output_MAC_6_32, output_MAC_6_33, output_MAC_6_34, output_MAC_6_35, output_MAC_6_36, output_MAC_6_37, output_MAC_6_38, output_MAC_6_39, 
		output_MAC_6_40, output_MAC_6_41, output_MAC_6_42, output_MAC_6_43, output_MAC_6_44, output_MAC_6_45, output_MAC_6_46, output_MAC_6_47, output_MAC_6_48, output_MAC_6_49, 
		output_MAC_6_50, output_MAC_6_51, output_MAC_6_52, output_MAC_6_53, output_MAC_6_54, output_MAC_6_55, output_MAC_6_56, output_MAC_6_57, output_MAC_6_58, output_MAC_6_59, 
		output_MAC_6_60, output_MAC_6_61, output_MAC_6_62, output_MAC_6_63, output_MAC_6_64, output_MAC_6_65, output_MAC_6_66, output_MAC_6_67, output_MAC_6_68, output_MAC_6_69, 
		output_MAC_6_70, output_MAC_6_71, output_MAC_6_72, output_MAC_6_73, output_MAC_6_74, output_MAC_6_75, output_MAC_6_76, output_MAC_6_77, output_MAC_6_78, output_MAC_6_79, 
		output_MAC_6_80, output_MAC_6_81, output_MAC_6_82, output_MAC_6_83, output_MAC_6_84, output_MAC_6_85, output_MAC_6_86, output_MAC_6_87, output_MAC_6_88, output_MAC_6_89, 
		output_MAC_6_90, output_MAC_6_91, output_MAC_6_92, output_MAC_6_93, output_MAC_6_94, output_MAC_6_95, output_MAC_6_96, output_MAC_6_97, output_MAC_6_98, output_MAC_6_99, 
		output_MAC_6_100, output_MAC_6_101, output_MAC_6_102, output_MAC_6_103, output_MAC_6_104, output_MAC_6_105, output_MAC_6_106, output_MAC_6_107, output_MAC_6_108, output_MAC_6_109, 
		output_MAC_6_110, output_MAC_6_111, output_MAC_6_112, output_MAC_6_113, output_MAC_6_114, output_MAC_6_115, output_MAC_6_116, output_MAC_6_117, output_MAC_6_118, output_MAC_6_119, 
		output_MAC_6_120, output_MAC_6_121, output_MAC_6_122, output_MAC_6_123, output_MAC_6_124, output_MAC_6_125, output_MAC_6_126, output_MAC_6_127, output_MAC_6_128, output_MAC_6_129, 
		output_MAC_6_130, output_MAC_6_131, output_MAC_6_132, output_MAC_6_133, output_MAC_6_134, output_MAC_6_135, output_MAC_6_136, output_MAC_6_137, output_MAC_6_138, output_MAC_6_139, 
		output_MAC_6_140, output_MAC_6_141, output_MAC_6_142, output_MAC_6_143, output_MAC_6_144, output_MAC_6_145, output_MAC_6_146, output_MAC_6_147, output_MAC_6_148, output_MAC_6_149, 
		output_MAC_6_150, output_MAC_6_151, output_MAC_6_152, output_MAC_6_153, output_MAC_6_154, output_MAC_6_155, output_MAC_6_156, output_MAC_6_157, output_MAC_6_158, output_MAC_6_159, 
		output_MAC_6_160, output_MAC_6_161, output_MAC_6_162, output_MAC_6_163, output_MAC_6_164, output_MAC_6_165, output_MAC_6_166, output_MAC_6_167, output_MAC_6_168, output_MAC_6_169, 
		output_MAC_6_170, output_MAC_6_171, output_MAC_6_172, output_MAC_6_173, output_MAC_6_174, output_MAC_6_175, output_MAC_6_176, output_MAC_6_177, output_MAC_6_178, output_MAC_6_179, 
		output_MAC_6_180, output_MAC_6_181, output_MAC_6_182, output_MAC_6_183, output_MAC_6_184, output_MAC_6_185, output_MAC_6_186, output_MAC_6_187, output_MAC_6_188, output_MAC_6_189, 
		output_MAC_6_190, output_MAC_6_191, output_MAC_6_192, output_MAC_6_193, output_MAC_6_194, output_MAC_6_195, output_MAC_6_196, output_MAC_6_197, output_MAC_6_198, output_MAC_6_199, 
		output_MAC_6_200, output_MAC_6_201, output_MAC_6_202, output_MAC_6_203, output_MAC_6_204, output_MAC_6_205, output_MAC_6_206, output_MAC_6_207, output_MAC_6_208, output_MAC_6_209, 
		output_MAC_6_210, output_MAC_6_211, output_MAC_6_212, output_MAC_6_213, output_MAC_6_214, output_MAC_6_215, output_MAC_6_216, output_MAC_6_217, output_MAC_6_218, output_MAC_6_219, 
		output_MAC_6_220, output_MAC_6_221, output_MAC_6_222, output_MAC_6_223, output_MAC_6_224, output_MAC_6_225, output_MAC_6_226, output_MAC_6_227, output_MAC_6_228, output_MAC_6_229, 
		output_MAC_6_230, output_MAC_6_231, output_MAC_6_232, output_MAC_6_233, output_MAC_6_234, output_MAC_6_235, output_MAC_6_236, output_MAC_6_237, output_MAC_6_238, output_MAC_6_239, 
		output_MAC_6_240, output_MAC_6_241, output_MAC_6_242, output_MAC_6_243, output_MAC_6_244, output_MAC_6_245, output_MAC_6_246, output_MAC_6_247, output_MAC_6_248, output_MAC_6_249, 
		output_MAC_6_250, output_MAC_6_251, output_MAC_6_252, output_MAC_6_253, output_MAC_6_254, output_MAC_6_255, output_MAC_6_256, output_MAC_6_257, output_MAC_6_258, output_MAC_6_259, 
		output_MAC_6_260, output_MAC_6_261, output_MAC_6_262, output_MAC_6_263, output_MAC_6_264, output_MAC_6_265, output_MAC_6_266, output_MAC_6_267, output_MAC_6_268, output_MAC_6_269, 
		output_MAC_6_270, output_MAC_6_271, output_MAC_6_272, output_MAC_6_273, output_MAC_6_274, output_MAC_6_275, output_MAC_6_276, output_MAC_6_277, output_MAC_6_278, output_MAC_6_279, 
		output_MAC_6_280, output_MAC_6_281, output_MAC_6_282, output_MAC_6_283, output_MAC_6_284, output_MAC_6_285, output_MAC_6_286, output_MAC_6_287, output_MAC_6_288, output_MAC_6_289, 
		output_MAC_6_290, output_MAC_6_291, output_MAC_6_292, output_MAC_6_293, output_MAC_6_294, output_MAC_6_295, output_MAC_6_296, output_MAC_6_297, output_MAC_6_298, output_MAC_6_299, 
		output_MAC_6_300, output_MAC_6_301, output_MAC_6_302, output_MAC_6_303, output_MAC_6_304, output_MAC_6_305, output_MAC_6_306, output_MAC_6_307, output_MAC_6_308, output_MAC_6_309, 
		output_MAC_6_310, output_MAC_6_311, output_MAC_6_312, output_MAC_6_313, output_MAC_6_314, output_MAC_6_315, output_MAC_6_316, output_MAC_6_317, output_MAC_6_318, output_MAC_6_319, 
		output_MAC_6_320, output_MAC_6_321, output_MAC_6_322, output_MAC_6_323, output_MAC_6_324, output_MAC_6_325, output_MAC_6_326, output_MAC_6_327, output_MAC_6_328, output_MAC_6_329, 
		output_MAC_6_330, output_MAC_6_331, output_MAC_6_332, output_MAC_6_333, output_MAC_6_334, output_MAC_6_335, output_MAC_6_336, output_MAC_6_337, output_MAC_6_338, output_MAC_6_339, 
		output_MAC_6_340, output_MAC_6_341, output_MAC_6_342, output_MAC_6_343, output_MAC_6_344, output_MAC_6_345, output_MAC_6_346, output_MAC_6_347, output_MAC_6_348, output_MAC_6_349, 
		output_MAC_6_350, output_MAC_6_351, output_MAC_6_352, output_MAC_6_353, output_MAC_6_354, output_MAC_6_355, output_MAC_6_356, output_MAC_6_357, output_MAC_6_358, output_MAC_6_359, 
		output_MAC_6_360, output_MAC_6_361, output_MAC_6_362, output_MAC_6_363, output_MAC_6_364, output_MAC_6_365, output_MAC_6_366, output_MAC_6_367, output_MAC_6_368, output_MAC_6_369, 
		output_MAC_6_370, output_MAC_6_371, output_MAC_6_372, output_MAC_6_373, output_MAC_6_374, output_MAC_6_375, output_MAC_6_376, output_MAC_6_377, output_MAC_6_378, output_MAC_6_379, 
		output_MAC_6_380, output_MAC_6_381, output_MAC_6_382, output_MAC_6_383, output_MAC_6_384, output_MAC_6_385, output_MAC_6_386, output_MAC_6_387, output_MAC_6_388, output_MAC_6_389, 
		output_MAC_6_390, output_MAC_6_391, output_MAC_6_392, output_MAC_6_393, output_MAC_6_394, output_MAC_6_395, output_MAC_6_396, output_MAC_6_397, output_MAC_6_398, output_MAC_6_399, 
		output_MAC_6_400, output_MAC_6_401, output_MAC_6_402, output_MAC_6_403, output_MAC_6_404, output_MAC_6_405, output_MAC_6_406, output_MAC_6_407, output_MAC_6_408, output_MAC_6_409, 
		output_MAC_6_410, output_MAC_6_411, output_MAC_6_412, output_MAC_6_413, output_MAC_6_414, output_MAC_6_415, output_MAC_6_416, output_MAC_6_417, output_MAC_6_418, output_MAC_6_419, 
		output_MAC_6_420, output_MAC_6_421, output_MAC_6_422, output_MAC_6_423, output_MAC_6_424, output_MAC_6_425, output_MAC_6_426, output_MAC_6_427, output_MAC_6_428, output_MAC_6_429, 
		output_MAC_6_430, output_MAC_6_431, output_MAC_6_432, output_MAC_6_433, output_MAC_6_434, output_MAC_6_435, output_MAC_6_436, output_MAC_6_437, output_MAC_6_438, output_MAC_6_439, 
		output_MAC_6_440, output_MAC_6_441, output_MAC_6_442, output_MAC_6_443, output_MAC_6_444, output_MAC_6_445, output_MAC_6_446, output_MAC_6_447, output_MAC_6_448, output_MAC_6_449, 
		output_MAC_6_450, output_MAC_6_451, output_MAC_6_452, output_MAC_6_453, output_MAC_6_454, output_MAC_6_455, output_MAC_6_456, output_MAC_6_457, output_MAC_6_458, output_MAC_6_459, 
		output_MAC_6_460, output_MAC_6_461, output_MAC_6_462, output_MAC_6_463, output_MAC_6_464, output_MAC_6_465, output_MAC_6_466, output_MAC_6_467, output_MAC_6_468, output_MAC_6_469, 
		output_MAC_6_470, output_MAC_6_471, output_MAC_6_472, output_MAC_6_473, output_MAC_6_474, output_MAC_6_475, output_MAC_6_476, output_MAC_6_477, output_MAC_6_478, output_MAC_6_479, 
		output_MAC_6_480, output_MAC_6_481, output_MAC_6_482, output_MAC_6_483, output_MAC_6_484, output_MAC_6_485, output_MAC_6_486, output_MAC_6_487, output_MAC_6_488, output_MAC_6_489, 
		output_MAC_6_490, output_MAC_6_491, output_MAC_6_492, output_MAC_6_493, output_MAC_6_494, output_MAC_6_495, output_MAC_6_496, output_MAC_6_497, output_MAC_6_498, output_MAC_6_499, 
		output_MAC_6_500, output_MAC_6_501, output_MAC_6_502, output_MAC_6_503, output_MAC_6_504, output_MAC_6_505, output_MAC_6_506, output_MAC_6_507, output_MAC_6_508, output_MAC_6_509, 
		output_MAC_6_510, output_MAC_6_511, output_MAC_6_512, output_MAC_6_513, output_MAC_6_514, output_MAC_6_515, output_MAC_6_516, output_MAC_6_517, output_MAC_6_518, output_MAC_6_519, 
		output_MAC_6_520, output_MAC_6_521, output_MAC_6_522, output_MAC_6_523, output_MAC_6_524, output_MAC_6_525, output_MAC_6_526, output_MAC_6_527, output_MAC_6_528, output_MAC_6_529, 
		output_MAC_6_530, output_MAC_6_531, output_MAC_6_532, output_MAC_6_533, output_MAC_6_534, output_MAC_6_535, output_MAC_6_536, output_MAC_6_537, output_MAC_6_538, output_MAC_6_539, 
		output_MAC_6_540, output_MAC_6_541, output_MAC_6_542, output_MAC_6_543, output_MAC_6_544, output_MAC_6_545, output_MAC_6_546, output_MAC_6_547, output_MAC_6_548, output_MAC_6_549, 
		output_MAC_6_550, output_MAC_6_551, output_MAC_6_552, output_MAC_6_553, output_MAC_6_554, output_MAC_6_555, output_MAC_6_556, output_MAC_6_557, output_MAC_6_558, output_MAC_6_559, 
		output_MAC_6_560, output_MAC_6_561, output_MAC_6_562, output_MAC_6_563, output_MAC_6_564, output_MAC_6_565, output_MAC_6_566, output_MAC_6_567, output_MAC_6_568, output_MAC_6_569, 
		output_MAC_6_570, output_MAC_6_571, output_MAC_6_572, output_MAC_6_573, output_MAC_6_574, output_MAC_6_575, output_MAC_6_576, output_MAC_6_577, output_MAC_6_578, output_MAC_6_579, 
		output_MAC_6_580, output_MAC_6_581, output_MAC_6_582, output_MAC_6_583, output_MAC_6_584, output_MAC_6_585, output_MAC_6_586, output_MAC_6_587, output_MAC_6_588, output_MAC_6_589, 
		output_MAC_6_590, output_MAC_6_591, output_MAC_6_592, output_MAC_6_593, output_MAC_6_594, output_MAC_6_595, output_MAC_6_596, output_MAC_6_597, output_MAC_6_598, output_MAC_6_599, 
		output_MAC_6_600, output_MAC_6_601, output_MAC_6_602, output_MAC_6_603, output_MAC_6_604, output_MAC_6_605, output_MAC_6_606, output_MAC_6_607, output_MAC_6_608, output_MAC_6_609, 
		output_MAC_6_610, output_MAC_6_611, output_MAC_6_612, output_MAC_6_613, output_MAC_6_614, output_MAC_6_615, output_MAC_6_616, output_MAC_6_617, output_MAC_6_618, output_MAC_6_619, 
		output_MAC_6_620, output_MAC_6_621, output_MAC_6_622, output_MAC_6_623, output_MAC_6_624, output_MAC_6_625, output_MAC_6_626, output_MAC_6_627, output_MAC_6_628, output_MAC_6_629, 
		output_MAC_6_630, output_MAC_6_631, output_MAC_6_632, output_MAC_6_633, output_MAC_6_634, output_MAC_6_635, output_MAC_6_636, output_MAC_6_637, output_MAC_6_638, output_MAC_6_639, 
		output_MAC_6_640, output_MAC_6_641, output_MAC_6_642, output_MAC_6_643, output_MAC_6_644, output_MAC_6_645, output_MAC_6_646, output_MAC_6_647, output_MAC_6_648, output_MAC_6_649, 
		output_MAC_6_650, output_MAC_6_651, output_MAC_6_652, output_MAC_6_653, output_MAC_6_654, output_MAC_6_655, output_MAC_6_656, output_MAC_6_657, output_MAC_6_658, output_MAC_6_659, 
		output_MAC_6_660, output_MAC_6_661, output_MAC_6_662, output_MAC_6_663, output_MAC_6_664, output_MAC_6_665, output_MAC_6_666, output_MAC_6_667, output_MAC_6_668, output_MAC_6_669, 
		output_MAC_6_670, output_MAC_6_671, output_MAC_6_672, output_MAC_6_673, output_MAC_6_674, output_MAC_6_675, output_MAC_6_676, output_MAC_6_677, output_MAC_6_678, output_MAC_6_679, 
		output_MAC_6_680, output_MAC_6_681, output_MAC_6_682, output_MAC_6_683, output_MAC_6_684, output_MAC_6_685, output_MAC_6_686, output_MAC_6_687, output_MAC_6_688, output_MAC_6_689, 
		output_MAC_6_690, output_MAC_6_691, output_MAC_6_692, output_MAC_6_693, output_MAC_6_694, output_MAC_6_695, output_MAC_6_696, output_MAC_6_697, output_MAC_6_698, output_MAC_6_699, 
		output_MAC_6_700, output_MAC_6_701, output_MAC_6_702, output_MAC_6_703, output_MAC_6_704, output_MAC_6_705, output_MAC_6_706, output_MAC_6_707, output_MAC_6_708, output_MAC_6_709, 
		output_MAC_6_710, output_MAC_6_711, output_MAC_6_712, output_MAC_6_713, output_MAC_6_714, output_MAC_6_715, output_MAC_6_716, output_MAC_6_717, output_MAC_6_718, output_MAC_6_719, 
		output_MAC_6_720, output_MAC_6_721, output_MAC_6_722, output_MAC_6_723, output_MAC_6_724, output_MAC_6_725, output_MAC_6_726, output_MAC_6_727, output_MAC_6_728, output_MAC_6_729, 
		output_MAC_6_730, output_MAC_6_731, output_MAC_6_732, output_MAC_6_733, output_MAC_6_734, output_MAC_6_735, output_MAC_6_736, output_MAC_6_737, output_MAC_6_738, output_MAC_6_739, 
		output_MAC_6_740, output_MAC_6_741, output_MAC_6_742, output_MAC_6_743, output_MAC_6_744, output_MAC_6_745, output_MAC_6_746, output_MAC_6_747, output_MAC_6_748, output_MAC_6_749, 
		output_MAC_6_750, output_MAC_6_751, output_MAC_6_752, output_MAC_6_753, output_MAC_6_754, output_MAC_6_755, output_MAC_6_756, output_MAC_6_757, output_MAC_6_758, output_MAC_6_759, 
		output_MAC_6_760, output_MAC_6_761, output_MAC_6_762, output_MAC_6_763, output_MAC_6_764, output_MAC_6_765, output_MAC_6_766, output_MAC_6_767: STD_LOGIC_VECTOR(31 downto 0);
	SIGNAL output_MAC_7_0, output_MAC_7_1, output_MAC_7_2, output_MAC_7_3, output_MAC_7_4, output_MAC_7_5, output_MAC_7_6, output_MAC_7_7, output_MAC_7_8, output_MAC_7_9, 
		output_MAC_7_10, output_MAC_7_11, output_MAC_7_12, output_MAC_7_13, output_MAC_7_14, output_MAC_7_15, output_MAC_7_16, output_MAC_7_17, output_MAC_7_18, output_MAC_7_19, 
		output_MAC_7_20, output_MAC_7_21, output_MAC_7_22, output_MAC_7_23, output_MAC_7_24, output_MAC_7_25, output_MAC_7_26, output_MAC_7_27, output_MAC_7_28, output_MAC_7_29, 
		output_MAC_7_30, output_MAC_7_31, output_MAC_7_32, output_MAC_7_33, output_MAC_7_34, output_MAC_7_35, output_MAC_7_36, output_MAC_7_37, output_MAC_7_38, output_MAC_7_39, 
		output_MAC_7_40, output_MAC_7_41, output_MAC_7_42, output_MAC_7_43, output_MAC_7_44, output_MAC_7_45, output_MAC_7_46, output_MAC_7_47, output_MAC_7_48, output_MAC_7_49, 
		output_MAC_7_50, output_MAC_7_51, output_MAC_7_52, output_MAC_7_53, output_MAC_7_54, output_MAC_7_55, output_MAC_7_56, output_MAC_7_57, output_MAC_7_58, output_MAC_7_59, 
		output_MAC_7_60, output_MAC_7_61, output_MAC_7_62, output_MAC_7_63, output_MAC_7_64, output_MAC_7_65, output_MAC_7_66, output_MAC_7_67, output_MAC_7_68, output_MAC_7_69, 
		output_MAC_7_70, output_MAC_7_71, output_MAC_7_72, output_MAC_7_73, output_MAC_7_74, output_MAC_7_75, output_MAC_7_76, output_MAC_7_77, output_MAC_7_78, output_MAC_7_79, 
		output_MAC_7_80, output_MAC_7_81, output_MAC_7_82, output_MAC_7_83, output_MAC_7_84, output_MAC_7_85, output_MAC_7_86, output_MAC_7_87, output_MAC_7_88, output_MAC_7_89, 
		output_MAC_7_90, output_MAC_7_91, output_MAC_7_92, output_MAC_7_93, output_MAC_7_94, output_MAC_7_95, output_MAC_7_96, output_MAC_7_97, output_MAC_7_98, output_MAC_7_99, 
		output_MAC_7_100, output_MAC_7_101, output_MAC_7_102, output_MAC_7_103, output_MAC_7_104, output_MAC_7_105, output_MAC_7_106, output_MAC_7_107, output_MAC_7_108, output_MAC_7_109, 
		output_MAC_7_110, output_MAC_7_111, output_MAC_7_112, output_MAC_7_113, output_MAC_7_114, output_MAC_7_115, output_MAC_7_116, output_MAC_7_117, output_MAC_7_118, output_MAC_7_119, 
		output_MAC_7_120, output_MAC_7_121, output_MAC_7_122, output_MAC_7_123, output_MAC_7_124, output_MAC_7_125, output_MAC_7_126, output_MAC_7_127, output_MAC_7_128, output_MAC_7_129, 
		output_MAC_7_130, output_MAC_7_131, output_MAC_7_132, output_MAC_7_133, output_MAC_7_134, output_MAC_7_135, output_MAC_7_136, output_MAC_7_137, output_MAC_7_138, output_MAC_7_139, 
		output_MAC_7_140, output_MAC_7_141, output_MAC_7_142, output_MAC_7_143, output_MAC_7_144, output_MAC_7_145, output_MAC_7_146, output_MAC_7_147, output_MAC_7_148, output_MAC_7_149, 
		output_MAC_7_150, output_MAC_7_151, output_MAC_7_152, output_MAC_7_153, output_MAC_7_154, output_MAC_7_155, output_MAC_7_156, output_MAC_7_157, output_MAC_7_158, output_MAC_7_159, 
		output_MAC_7_160, output_MAC_7_161, output_MAC_7_162, output_MAC_7_163, output_MAC_7_164, output_MAC_7_165, output_MAC_7_166, output_MAC_7_167, output_MAC_7_168, output_MAC_7_169, 
		output_MAC_7_170, output_MAC_7_171, output_MAC_7_172, output_MAC_7_173, output_MAC_7_174, output_MAC_7_175, output_MAC_7_176, output_MAC_7_177, output_MAC_7_178, output_MAC_7_179, 
		output_MAC_7_180, output_MAC_7_181, output_MAC_7_182, output_MAC_7_183, output_MAC_7_184, output_MAC_7_185, output_MAC_7_186, output_MAC_7_187, output_MAC_7_188, output_MAC_7_189, 
		output_MAC_7_190, output_MAC_7_191, output_MAC_7_192, output_MAC_7_193, output_MAC_7_194, output_MAC_7_195, output_MAC_7_196, output_MAC_7_197, output_MAC_7_198, output_MAC_7_199, 
		output_MAC_7_200, output_MAC_7_201, output_MAC_7_202, output_MAC_7_203, output_MAC_7_204, output_MAC_7_205, output_MAC_7_206, output_MAC_7_207, output_MAC_7_208, output_MAC_7_209, 
		output_MAC_7_210, output_MAC_7_211, output_MAC_7_212, output_MAC_7_213, output_MAC_7_214, output_MAC_7_215, output_MAC_7_216, output_MAC_7_217, output_MAC_7_218, output_MAC_7_219, 
		output_MAC_7_220, output_MAC_7_221, output_MAC_7_222, output_MAC_7_223, output_MAC_7_224, output_MAC_7_225, output_MAC_7_226, output_MAC_7_227, output_MAC_7_228, output_MAC_7_229, 
		output_MAC_7_230, output_MAC_7_231, output_MAC_7_232, output_MAC_7_233, output_MAC_7_234, output_MAC_7_235, output_MAC_7_236, output_MAC_7_237, output_MAC_7_238, output_MAC_7_239, 
		output_MAC_7_240, output_MAC_7_241, output_MAC_7_242, output_MAC_7_243, output_MAC_7_244, output_MAC_7_245, output_MAC_7_246, output_MAC_7_247, output_MAC_7_248, output_MAC_7_249, 
		output_MAC_7_250, output_MAC_7_251, output_MAC_7_252, output_MAC_7_253, output_MAC_7_254, output_MAC_7_255, output_MAC_7_256, output_MAC_7_257, output_MAC_7_258, output_MAC_7_259, 
		output_MAC_7_260, output_MAC_7_261, output_MAC_7_262, output_MAC_7_263, output_MAC_7_264, output_MAC_7_265, output_MAC_7_266, output_MAC_7_267, output_MAC_7_268, output_MAC_7_269, 
		output_MAC_7_270, output_MAC_7_271, output_MAC_7_272, output_MAC_7_273, output_MAC_7_274, output_MAC_7_275, output_MAC_7_276, output_MAC_7_277, output_MAC_7_278, output_MAC_7_279, 
		output_MAC_7_280, output_MAC_7_281, output_MAC_7_282, output_MAC_7_283, output_MAC_7_284, output_MAC_7_285, output_MAC_7_286, output_MAC_7_287, output_MAC_7_288, output_MAC_7_289, 
		output_MAC_7_290, output_MAC_7_291, output_MAC_7_292, output_MAC_7_293, output_MAC_7_294, output_MAC_7_295, output_MAC_7_296, output_MAC_7_297, output_MAC_7_298, output_MAC_7_299, 
		output_MAC_7_300, output_MAC_7_301, output_MAC_7_302, output_MAC_7_303, output_MAC_7_304, output_MAC_7_305, output_MAC_7_306, output_MAC_7_307, output_MAC_7_308, output_MAC_7_309, 
		output_MAC_7_310, output_MAC_7_311, output_MAC_7_312, output_MAC_7_313, output_MAC_7_314, output_MAC_7_315, output_MAC_7_316, output_MAC_7_317, output_MAC_7_318, output_MAC_7_319, 
		output_MAC_7_320, output_MAC_7_321, output_MAC_7_322, output_MAC_7_323, output_MAC_7_324, output_MAC_7_325, output_MAC_7_326, output_MAC_7_327, output_MAC_7_328, output_MAC_7_329, 
		output_MAC_7_330, output_MAC_7_331, output_MAC_7_332, output_MAC_7_333, output_MAC_7_334, output_MAC_7_335, output_MAC_7_336, output_MAC_7_337, output_MAC_7_338, output_MAC_7_339, 
		output_MAC_7_340, output_MAC_7_341, output_MAC_7_342, output_MAC_7_343, output_MAC_7_344, output_MAC_7_345, output_MAC_7_346, output_MAC_7_347, output_MAC_7_348, output_MAC_7_349, 
		output_MAC_7_350, output_MAC_7_351, output_MAC_7_352, output_MAC_7_353, output_MAC_7_354, output_MAC_7_355, output_MAC_7_356, output_MAC_7_357, output_MAC_7_358, output_MAC_7_359, 
		output_MAC_7_360, output_MAC_7_361, output_MAC_7_362, output_MAC_7_363, output_MAC_7_364, output_MAC_7_365, output_MAC_7_366, output_MAC_7_367, output_MAC_7_368, output_MAC_7_369, 
		output_MAC_7_370, output_MAC_7_371, output_MAC_7_372, output_MAC_7_373, output_MAC_7_374, output_MAC_7_375, output_MAC_7_376, output_MAC_7_377, output_MAC_7_378, output_MAC_7_379, 
		output_MAC_7_380, output_MAC_7_381, output_MAC_7_382, output_MAC_7_383, output_MAC_7_384, output_MAC_7_385, output_MAC_7_386, output_MAC_7_387, output_MAC_7_388, output_MAC_7_389, 
		output_MAC_7_390, output_MAC_7_391, output_MAC_7_392, output_MAC_7_393, output_MAC_7_394, output_MAC_7_395, output_MAC_7_396, output_MAC_7_397, output_MAC_7_398, output_MAC_7_399, 
		output_MAC_7_400, output_MAC_7_401, output_MAC_7_402, output_MAC_7_403, output_MAC_7_404, output_MAC_7_405, output_MAC_7_406, output_MAC_7_407, output_MAC_7_408, output_MAC_7_409, 
		output_MAC_7_410, output_MAC_7_411, output_MAC_7_412, output_MAC_7_413, output_MAC_7_414, output_MAC_7_415, output_MAC_7_416, output_MAC_7_417, output_MAC_7_418, output_MAC_7_419, 
		output_MAC_7_420, output_MAC_7_421, output_MAC_7_422, output_MAC_7_423, output_MAC_7_424, output_MAC_7_425, output_MAC_7_426, output_MAC_7_427, output_MAC_7_428, output_MAC_7_429, 
		output_MAC_7_430, output_MAC_7_431, output_MAC_7_432, output_MAC_7_433, output_MAC_7_434, output_MAC_7_435, output_MAC_7_436, output_MAC_7_437, output_MAC_7_438, output_MAC_7_439, 
		output_MAC_7_440, output_MAC_7_441, output_MAC_7_442, output_MAC_7_443, output_MAC_7_444, output_MAC_7_445, output_MAC_7_446, output_MAC_7_447, output_MAC_7_448, output_MAC_7_449, 
		output_MAC_7_450, output_MAC_7_451, output_MAC_7_452, output_MAC_7_453, output_MAC_7_454, output_MAC_7_455, output_MAC_7_456, output_MAC_7_457, output_MAC_7_458, output_MAC_7_459, 
		output_MAC_7_460, output_MAC_7_461, output_MAC_7_462, output_MAC_7_463, output_MAC_7_464, output_MAC_7_465, output_MAC_7_466, output_MAC_7_467, output_MAC_7_468, output_MAC_7_469, 
		output_MAC_7_470, output_MAC_7_471, output_MAC_7_472, output_MAC_7_473, output_MAC_7_474, output_MAC_7_475, output_MAC_7_476, output_MAC_7_477, output_MAC_7_478, output_MAC_7_479, 
		output_MAC_7_480, output_MAC_7_481, output_MAC_7_482, output_MAC_7_483, output_MAC_7_484, output_MAC_7_485, output_MAC_7_486, output_MAC_7_487, output_MAC_7_488, output_MAC_7_489, 
		output_MAC_7_490, output_MAC_7_491, output_MAC_7_492, output_MAC_7_493, output_MAC_7_494, output_MAC_7_495, output_MAC_7_496, output_MAC_7_497, output_MAC_7_498, output_MAC_7_499, 
		output_MAC_7_500, output_MAC_7_501, output_MAC_7_502, output_MAC_7_503, output_MAC_7_504, output_MAC_7_505, output_MAC_7_506, output_MAC_7_507, output_MAC_7_508, output_MAC_7_509, 
		output_MAC_7_510, output_MAC_7_511, output_MAC_7_512, output_MAC_7_513, output_MAC_7_514, output_MAC_7_515, output_MAC_7_516, output_MAC_7_517, output_MAC_7_518, output_MAC_7_519, 
		output_MAC_7_520, output_MAC_7_521, output_MAC_7_522, output_MAC_7_523, output_MAC_7_524, output_MAC_7_525, output_MAC_7_526, output_MAC_7_527, output_MAC_7_528, output_MAC_7_529, 
		output_MAC_7_530, output_MAC_7_531, output_MAC_7_532, output_MAC_7_533, output_MAC_7_534, output_MAC_7_535, output_MAC_7_536, output_MAC_7_537, output_MAC_7_538, output_MAC_7_539, 
		output_MAC_7_540, output_MAC_7_541, output_MAC_7_542, output_MAC_7_543, output_MAC_7_544, output_MAC_7_545, output_MAC_7_546, output_MAC_7_547, output_MAC_7_548, output_MAC_7_549, 
		output_MAC_7_550, output_MAC_7_551, output_MAC_7_552, output_MAC_7_553, output_MAC_7_554, output_MAC_7_555, output_MAC_7_556, output_MAC_7_557, output_MAC_7_558, output_MAC_7_559, 
		output_MAC_7_560, output_MAC_7_561, output_MAC_7_562, output_MAC_7_563, output_MAC_7_564, output_MAC_7_565, output_MAC_7_566, output_MAC_7_567, output_MAC_7_568, output_MAC_7_569, 
		output_MAC_7_570, output_MAC_7_571, output_MAC_7_572, output_MAC_7_573, output_MAC_7_574, output_MAC_7_575, output_MAC_7_576, output_MAC_7_577, output_MAC_7_578, output_MAC_7_579, 
		output_MAC_7_580, output_MAC_7_581, output_MAC_7_582, output_MAC_7_583, output_MAC_7_584, output_MAC_7_585, output_MAC_7_586, output_MAC_7_587, output_MAC_7_588, output_MAC_7_589, 
		output_MAC_7_590, output_MAC_7_591, output_MAC_7_592, output_MAC_7_593, output_MAC_7_594, output_MAC_7_595, output_MAC_7_596, output_MAC_7_597, output_MAC_7_598, output_MAC_7_599, 
		output_MAC_7_600, output_MAC_7_601, output_MAC_7_602, output_MAC_7_603, output_MAC_7_604, output_MAC_7_605, output_MAC_7_606, output_MAC_7_607, output_MAC_7_608, output_MAC_7_609, 
		output_MAC_7_610, output_MAC_7_611, output_MAC_7_612, output_MAC_7_613, output_MAC_7_614, output_MAC_7_615, output_MAC_7_616, output_MAC_7_617, output_MAC_7_618, output_MAC_7_619, 
		output_MAC_7_620, output_MAC_7_621, output_MAC_7_622, output_MAC_7_623, output_MAC_7_624, output_MAC_7_625, output_MAC_7_626, output_MAC_7_627, output_MAC_7_628, output_MAC_7_629, 
		output_MAC_7_630, output_MAC_7_631, output_MAC_7_632, output_MAC_7_633, output_MAC_7_634, output_MAC_7_635, output_MAC_7_636, output_MAC_7_637, output_MAC_7_638, output_MAC_7_639, 
		output_MAC_7_640, output_MAC_7_641, output_MAC_7_642, output_MAC_7_643, output_MAC_7_644, output_MAC_7_645, output_MAC_7_646, output_MAC_7_647, output_MAC_7_648, output_MAC_7_649, 
		output_MAC_7_650, output_MAC_7_651, output_MAC_7_652, output_MAC_7_653, output_MAC_7_654, output_MAC_7_655, output_MAC_7_656, output_MAC_7_657, output_MAC_7_658, output_MAC_7_659, 
		output_MAC_7_660, output_MAC_7_661, output_MAC_7_662, output_MAC_7_663, output_MAC_7_664, output_MAC_7_665, output_MAC_7_666, output_MAC_7_667, output_MAC_7_668, output_MAC_7_669, 
		output_MAC_7_670, output_MAC_7_671, output_MAC_7_672, output_MAC_7_673, output_MAC_7_674, output_MAC_7_675, output_MAC_7_676, output_MAC_7_677, output_MAC_7_678, output_MAC_7_679, 
		output_MAC_7_680, output_MAC_7_681, output_MAC_7_682, output_MAC_7_683, output_MAC_7_684, output_MAC_7_685, output_MAC_7_686, output_MAC_7_687, output_MAC_7_688, output_MAC_7_689, 
		output_MAC_7_690, output_MAC_7_691, output_MAC_7_692, output_MAC_7_693, output_MAC_7_694, output_MAC_7_695, output_MAC_7_696, output_MAC_7_697, output_MAC_7_698, output_MAC_7_699, 
		output_MAC_7_700, output_MAC_7_701, output_MAC_7_702, output_MAC_7_703, output_MAC_7_704, output_MAC_7_705, output_MAC_7_706, output_MAC_7_707, output_MAC_7_708, output_MAC_7_709, 
		output_MAC_7_710, output_MAC_7_711, output_MAC_7_712, output_MAC_7_713, output_MAC_7_714, output_MAC_7_715, output_MAC_7_716, output_MAC_7_717, output_MAC_7_718, output_MAC_7_719, 
		output_MAC_7_720, output_MAC_7_721, output_MAC_7_722, output_MAC_7_723, output_MAC_7_724, output_MAC_7_725, output_MAC_7_726, output_MAC_7_727, output_MAC_7_728, output_MAC_7_729, 
		output_MAC_7_730, output_MAC_7_731, output_MAC_7_732, output_MAC_7_733, output_MAC_7_734, output_MAC_7_735, output_MAC_7_736, output_MAC_7_737, output_MAC_7_738, output_MAC_7_739, 
		output_MAC_7_740, output_MAC_7_741, output_MAC_7_742, output_MAC_7_743, output_MAC_7_744, output_MAC_7_745, output_MAC_7_746, output_MAC_7_747, output_MAC_7_748, output_MAC_7_749, 
		output_MAC_7_750, output_MAC_7_751, output_MAC_7_752, output_MAC_7_753, output_MAC_7_754, output_MAC_7_755, output_MAC_7_756, output_MAC_7_757, output_MAC_7_758, output_MAC_7_759, 
		output_MAC_7_760, output_MAC_7_761, output_MAC_7_762, output_MAC_7_763, output_MAC_7_764, output_MAC_7_765, output_MAC_7_766, output_MAC_7_767: STD_LOGIC_VECTOR(31 downto 0);

BEGIN

	MAC_0_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_0, data_out=>output_MAC_0_0);
	MAC_0_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_1, data_out=>output_MAC_0_1);
	MAC_0_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_2, data_out=>output_MAC_0_2);
	MAC_0_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_3, data_out=>output_MAC_0_3);
	MAC_0_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_4, data_out=>output_MAC_0_4);
	MAC_0_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_5, data_out=>output_MAC_0_5);
	MAC_0_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_6, data_out=>output_MAC_0_6);
	MAC_0_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_7, data_out=>output_MAC_0_7);
	MAC_0_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_8, data_out=>output_MAC_0_8);
	MAC_0_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_9, data_out=>output_MAC_0_9);
	MAC_0_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_10, data_out=>output_MAC_0_10);
	MAC_0_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_11, data_out=>output_MAC_0_11);
	MAC_0_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_12, data_out=>output_MAC_0_12);
	MAC_0_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_13, data_out=>output_MAC_0_13);
	MAC_0_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_14, data_out=>output_MAC_0_14);
	MAC_0_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_15, data_out=>output_MAC_0_15);
	MAC_0_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_16, data_out=>output_MAC_0_16);
	MAC_0_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_17, data_out=>output_MAC_0_17);
	MAC_0_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_18, data_out=>output_MAC_0_18);
	MAC_0_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_19, data_out=>output_MAC_0_19);
	MAC_0_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_20, data_out=>output_MAC_0_20);
	MAC_0_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_21, data_out=>output_MAC_0_21);
	MAC_0_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_22, data_out=>output_MAC_0_22);
	MAC_0_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_23, data_out=>output_MAC_0_23);
	MAC_0_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_24, data_out=>output_MAC_0_24);
	MAC_0_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_25, data_out=>output_MAC_0_25);
	MAC_0_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_26, data_out=>output_MAC_0_26);
	MAC_0_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_27, data_out=>output_MAC_0_27);
	MAC_0_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_28, data_out=>output_MAC_0_28);
	MAC_0_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_29, data_out=>output_MAC_0_29);
	MAC_0_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_30, data_out=>output_MAC_0_30);
	MAC_0_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_31, data_out=>output_MAC_0_31);
	MAC_0_32: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_32, data_out=>output_MAC_0_32);
	MAC_0_33: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_33, data_out=>output_MAC_0_33);
	MAC_0_34: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_34, data_out=>output_MAC_0_34);
	MAC_0_35: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_35, data_out=>output_MAC_0_35);
	MAC_0_36: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_36, data_out=>output_MAC_0_36);
	MAC_0_37: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_37, data_out=>output_MAC_0_37);
	MAC_0_38: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_38, data_out=>output_MAC_0_38);
	MAC_0_39: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_39, data_out=>output_MAC_0_39);
	MAC_0_40: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_40, data_out=>output_MAC_0_40);
	MAC_0_41: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_41, data_out=>output_MAC_0_41);
	MAC_0_42: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_42, data_out=>output_MAC_0_42);
	MAC_0_43: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_43, data_out=>output_MAC_0_43);
	MAC_0_44: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_44, data_out=>output_MAC_0_44);
	MAC_0_45: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_45, data_out=>output_MAC_0_45);
	MAC_0_46: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_46, data_out=>output_MAC_0_46);
	MAC_0_47: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_47, data_out=>output_MAC_0_47);
	MAC_0_48: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_48, data_out=>output_MAC_0_48);
	MAC_0_49: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_49, data_out=>output_MAC_0_49);
	MAC_0_50: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_50, data_out=>output_MAC_0_50);
	MAC_0_51: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_51, data_out=>output_MAC_0_51);
	MAC_0_52: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_52, data_out=>output_MAC_0_52);
	MAC_0_53: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_53, data_out=>output_MAC_0_53);
	MAC_0_54: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_54, data_out=>output_MAC_0_54);
	MAC_0_55: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_55, data_out=>output_MAC_0_55);
	MAC_0_56: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_56, data_out=>output_MAC_0_56);
	MAC_0_57: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_57, data_out=>output_MAC_0_57);
	MAC_0_58: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_58, data_out=>output_MAC_0_58);
	MAC_0_59: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_59, data_out=>output_MAC_0_59);
	MAC_0_60: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_60, data_out=>output_MAC_0_60);
	MAC_0_61: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_61, data_out=>output_MAC_0_61);
	MAC_0_62: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_62, data_out=>output_MAC_0_62);
	MAC_0_63: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_63, data_out=>output_MAC_0_63);
	MAC_0_64: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_64, data_out=>output_MAC_0_64);
	MAC_0_65: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_65, data_out=>output_MAC_0_65);
	MAC_0_66: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_66, data_out=>output_MAC_0_66);
	MAC_0_67: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_67, data_out=>output_MAC_0_67);
	MAC_0_68: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_68, data_out=>output_MAC_0_68);
	MAC_0_69: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_69, data_out=>output_MAC_0_69);
	MAC_0_70: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_70, data_out=>output_MAC_0_70);
	MAC_0_71: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_71, data_out=>output_MAC_0_71);
	MAC_0_72: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_72, data_out=>output_MAC_0_72);
	MAC_0_73: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_73, data_out=>output_MAC_0_73);
	MAC_0_74: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_74, data_out=>output_MAC_0_74);
	MAC_0_75: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_75, data_out=>output_MAC_0_75);
	MAC_0_76: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_76, data_out=>output_MAC_0_76);
	MAC_0_77: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_77, data_out=>output_MAC_0_77);
	MAC_0_78: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_78, data_out=>output_MAC_0_78);
	MAC_0_79: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_79, data_out=>output_MAC_0_79);
	MAC_0_80: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_80, data_out=>output_MAC_0_80);
	MAC_0_81: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_81, data_out=>output_MAC_0_81);
	MAC_0_82: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_82, data_out=>output_MAC_0_82);
	MAC_0_83: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_83, data_out=>output_MAC_0_83);
	MAC_0_84: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_84, data_out=>output_MAC_0_84);
	MAC_0_85: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_85, data_out=>output_MAC_0_85);
	MAC_0_86: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_86, data_out=>output_MAC_0_86);
	MAC_0_87: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_87, data_out=>output_MAC_0_87);
	MAC_0_88: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_88, data_out=>output_MAC_0_88);
	MAC_0_89: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_89, data_out=>output_MAC_0_89);
	MAC_0_90: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_90, data_out=>output_MAC_0_90);
	MAC_0_91: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_91, data_out=>output_MAC_0_91);
	MAC_0_92: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_92, data_out=>output_MAC_0_92);
	MAC_0_93: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_93, data_out=>output_MAC_0_93);
	MAC_0_94: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_94, data_out=>output_MAC_0_94);
	MAC_0_95: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_95, data_out=>output_MAC_0_95);
	MAC_0_96: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_96, data_out=>output_MAC_0_96);
	MAC_0_97: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_97, data_out=>output_MAC_0_97);
	MAC_0_98: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_98, data_out=>output_MAC_0_98);
	MAC_0_99: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_99, data_out=>output_MAC_0_99);
	MAC_0_100: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_100, data_out=>output_MAC_0_100);
	MAC_0_101: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_101, data_out=>output_MAC_0_101);
	MAC_0_102: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_102, data_out=>output_MAC_0_102);
	MAC_0_103: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_103, data_out=>output_MAC_0_103);
	MAC_0_104: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_104, data_out=>output_MAC_0_104);
	MAC_0_105: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_105, data_out=>output_MAC_0_105);
	MAC_0_106: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_106, data_out=>output_MAC_0_106);
	MAC_0_107: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_107, data_out=>output_MAC_0_107);
	MAC_0_108: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_108, data_out=>output_MAC_0_108);
	MAC_0_109: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_109, data_out=>output_MAC_0_109);
	MAC_0_110: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_110, data_out=>output_MAC_0_110);
	MAC_0_111: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_111, data_out=>output_MAC_0_111);
	MAC_0_112: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_112, data_out=>output_MAC_0_112);
	MAC_0_113: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_113, data_out=>output_MAC_0_113);
	MAC_0_114: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_114, data_out=>output_MAC_0_114);
	MAC_0_115: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_115, data_out=>output_MAC_0_115);
	MAC_0_116: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_116, data_out=>output_MAC_0_116);
	MAC_0_117: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_117, data_out=>output_MAC_0_117);
	MAC_0_118: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_118, data_out=>output_MAC_0_118);
	MAC_0_119: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_119, data_out=>output_MAC_0_119);
	MAC_0_120: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_120, data_out=>output_MAC_0_120);
	MAC_0_121: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_121, data_out=>output_MAC_0_121);
	MAC_0_122: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_122, data_out=>output_MAC_0_122);
	MAC_0_123: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_123, data_out=>output_MAC_0_123);
	MAC_0_124: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_124, data_out=>output_MAC_0_124);
	MAC_0_125: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_125, data_out=>output_MAC_0_125);
	MAC_0_126: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_126, data_out=>output_MAC_0_126);
	MAC_0_127: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_127, data_out=>output_MAC_0_127);
	MAC_0_128: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_128, data_out=>output_MAC_0_128);
	MAC_0_129: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_129, data_out=>output_MAC_0_129);
	MAC_0_130: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_130, data_out=>output_MAC_0_130);
	MAC_0_131: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_131, data_out=>output_MAC_0_131);
	MAC_0_132: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_132, data_out=>output_MAC_0_132);
	MAC_0_133: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_133, data_out=>output_MAC_0_133);
	MAC_0_134: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_134, data_out=>output_MAC_0_134);
	MAC_0_135: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_135, data_out=>output_MAC_0_135);
	MAC_0_136: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_136, data_out=>output_MAC_0_136);
	MAC_0_137: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_137, data_out=>output_MAC_0_137);
	MAC_0_138: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_138, data_out=>output_MAC_0_138);
	MAC_0_139: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_139, data_out=>output_MAC_0_139);
	MAC_0_140: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_140, data_out=>output_MAC_0_140);
	MAC_0_141: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_141, data_out=>output_MAC_0_141);
	MAC_0_142: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_142, data_out=>output_MAC_0_142);
	MAC_0_143: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_143, data_out=>output_MAC_0_143);
	MAC_0_144: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_144, data_out=>output_MAC_0_144);
	MAC_0_145: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_145, data_out=>output_MAC_0_145);
	MAC_0_146: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_146, data_out=>output_MAC_0_146);
	MAC_0_147: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_147, data_out=>output_MAC_0_147);
	MAC_0_148: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_148, data_out=>output_MAC_0_148);
	MAC_0_149: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_149, data_out=>output_MAC_0_149);
	MAC_0_150: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_150, data_out=>output_MAC_0_150);
	MAC_0_151: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_151, data_out=>output_MAC_0_151);
	MAC_0_152: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_152, data_out=>output_MAC_0_152);
	MAC_0_153: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_153, data_out=>output_MAC_0_153);
	MAC_0_154: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_154, data_out=>output_MAC_0_154);
	MAC_0_155: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_155, data_out=>output_MAC_0_155);
	MAC_0_156: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_156, data_out=>output_MAC_0_156);
	MAC_0_157: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_157, data_out=>output_MAC_0_157);
	MAC_0_158: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_158, data_out=>output_MAC_0_158);
	MAC_0_159: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_159, data_out=>output_MAC_0_159);
	MAC_0_160: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_160, data_out=>output_MAC_0_160);
	MAC_0_161: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_161, data_out=>output_MAC_0_161);
	MAC_0_162: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_162, data_out=>output_MAC_0_162);
	MAC_0_163: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_163, data_out=>output_MAC_0_163);
	MAC_0_164: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_164, data_out=>output_MAC_0_164);
	MAC_0_165: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_165, data_out=>output_MAC_0_165);
	MAC_0_166: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_166, data_out=>output_MAC_0_166);
	MAC_0_167: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_167, data_out=>output_MAC_0_167);
	MAC_0_168: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_168, data_out=>output_MAC_0_168);
	MAC_0_169: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_169, data_out=>output_MAC_0_169);
	MAC_0_170: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_170, data_out=>output_MAC_0_170);
	MAC_0_171: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_171, data_out=>output_MAC_0_171);
	MAC_0_172: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_172, data_out=>output_MAC_0_172);
	MAC_0_173: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_173, data_out=>output_MAC_0_173);
	MAC_0_174: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_174, data_out=>output_MAC_0_174);
	MAC_0_175: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_175, data_out=>output_MAC_0_175);
	MAC_0_176: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_176, data_out=>output_MAC_0_176);
	MAC_0_177: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_177, data_out=>output_MAC_0_177);
	MAC_0_178: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_178, data_out=>output_MAC_0_178);
	MAC_0_179: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_179, data_out=>output_MAC_0_179);
	MAC_0_180: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_180, data_out=>output_MAC_0_180);
	MAC_0_181: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_181, data_out=>output_MAC_0_181);
	MAC_0_182: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_182, data_out=>output_MAC_0_182);
	MAC_0_183: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_183, data_out=>output_MAC_0_183);
	MAC_0_184: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_184, data_out=>output_MAC_0_184);
	MAC_0_185: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_185, data_out=>output_MAC_0_185);
	MAC_0_186: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_186, data_out=>output_MAC_0_186);
	MAC_0_187: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_187, data_out=>output_MAC_0_187);
	MAC_0_188: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_188, data_out=>output_MAC_0_188);
	MAC_0_189: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_189, data_out=>output_MAC_0_189);
	MAC_0_190: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_190, data_out=>output_MAC_0_190);
	MAC_0_191: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_191, data_out=>output_MAC_0_191);
	MAC_0_192: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_192, data_out=>output_MAC_0_192);
	MAC_0_193: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_193, data_out=>output_MAC_0_193);
	MAC_0_194: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_194, data_out=>output_MAC_0_194);
	MAC_0_195: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_195, data_out=>output_MAC_0_195);
	MAC_0_196: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_196, data_out=>output_MAC_0_196);
	MAC_0_197: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_197, data_out=>output_MAC_0_197);
	MAC_0_198: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_198, data_out=>output_MAC_0_198);
	MAC_0_199: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_199, data_out=>output_MAC_0_199);
	MAC_0_200: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_200, data_out=>output_MAC_0_200);
	MAC_0_201: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_201, data_out=>output_MAC_0_201);
	MAC_0_202: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_202, data_out=>output_MAC_0_202);
	MAC_0_203: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_203, data_out=>output_MAC_0_203);
	MAC_0_204: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_204, data_out=>output_MAC_0_204);
	MAC_0_205: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_205, data_out=>output_MAC_0_205);
	MAC_0_206: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_206, data_out=>output_MAC_0_206);
	MAC_0_207: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_207, data_out=>output_MAC_0_207);
	MAC_0_208: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_208, data_out=>output_MAC_0_208);
	MAC_0_209: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_209, data_out=>output_MAC_0_209);
	MAC_0_210: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_210, data_out=>output_MAC_0_210);
	MAC_0_211: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_211, data_out=>output_MAC_0_211);
	MAC_0_212: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_212, data_out=>output_MAC_0_212);
	MAC_0_213: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_213, data_out=>output_MAC_0_213);
	MAC_0_214: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_214, data_out=>output_MAC_0_214);
	MAC_0_215: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_215, data_out=>output_MAC_0_215);
	MAC_0_216: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_216, data_out=>output_MAC_0_216);
	MAC_0_217: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_217, data_out=>output_MAC_0_217);
	MAC_0_218: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_218, data_out=>output_MAC_0_218);
	MAC_0_219: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_219, data_out=>output_MAC_0_219);
	MAC_0_220: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_220, data_out=>output_MAC_0_220);
	MAC_0_221: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_221, data_out=>output_MAC_0_221);
	MAC_0_222: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_222, data_out=>output_MAC_0_222);
	MAC_0_223: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_223, data_out=>output_MAC_0_223);
	MAC_0_224: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_224, data_out=>output_MAC_0_224);
	MAC_0_225: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_225, data_out=>output_MAC_0_225);
	MAC_0_226: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_226, data_out=>output_MAC_0_226);
	MAC_0_227: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_227, data_out=>output_MAC_0_227);
	MAC_0_228: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_228, data_out=>output_MAC_0_228);
	MAC_0_229: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_229, data_out=>output_MAC_0_229);
	MAC_0_230: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_230, data_out=>output_MAC_0_230);
	MAC_0_231: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_231, data_out=>output_MAC_0_231);
	MAC_0_232: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_232, data_out=>output_MAC_0_232);
	MAC_0_233: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_233, data_out=>output_MAC_0_233);
	MAC_0_234: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_234, data_out=>output_MAC_0_234);
	MAC_0_235: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_235, data_out=>output_MAC_0_235);
	MAC_0_236: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_236, data_out=>output_MAC_0_236);
	MAC_0_237: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_237, data_out=>output_MAC_0_237);
	MAC_0_238: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_238, data_out=>output_MAC_0_238);
	MAC_0_239: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_239, data_out=>output_MAC_0_239);
	MAC_0_240: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_240, data_out=>output_MAC_0_240);
	MAC_0_241: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_241, data_out=>output_MAC_0_241);
	MAC_0_242: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_242, data_out=>output_MAC_0_242);
	MAC_0_243: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_243, data_out=>output_MAC_0_243);
	MAC_0_244: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_244, data_out=>output_MAC_0_244);
	MAC_0_245: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_245, data_out=>output_MAC_0_245);
	MAC_0_246: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_246, data_out=>output_MAC_0_246);
	MAC_0_247: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_247, data_out=>output_MAC_0_247);
	MAC_0_248: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_248, data_out=>output_MAC_0_248);
	MAC_0_249: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_249, data_out=>output_MAC_0_249);
	MAC_0_250: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_250, data_out=>output_MAC_0_250);
	MAC_0_251: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_251, data_out=>output_MAC_0_251);
	MAC_0_252: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_252, data_out=>output_MAC_0_252);
	MAC_0_253: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_253, data_out=>output_MAC_0_253);
	MAC_0_254: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_254, data_out=>output_MAC_0_254);
	MAC_0_255: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_255, data_out=>output_MAC_0_255);
	MAC_0_256: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_256, data_out=>output_MAC_0_256);
	MAC_0_257: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_257, data_out=>output_MAC_0_257);
	MAC_0_258: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_258, data_out=>output_MAC_0_258);
	MAC_0_259: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_259, data_out=>output_MAC_0_259);
	MAC_0_260: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_260, data_out=>output_MAC_0_260);
	MAC_0_261: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_261, data_out=>output_MAC_0_261);
	MAC_0_262: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_262, data_out=>output_MAC_0_262);
	MAC_0_263: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_263, data_out=>output_MAC_0_263);
	MAC_0_264: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_264, data_out=>output_MAC_0_264);
	MAC_0_265: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_265, data_out=>output_MAC_0_265);
	MAC_0_266: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_266, data_out=>output_MAC_0_266);
	MAC_0_267: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_267, data_out=>output_MAC_0_267);
	MAC_0_268: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_268, data_out=>output_MAC_0_268);
	MAC_0_269: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_269, data_out=>output_MAC_0_269);
	MAC_0_270: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_270, data_out=>output_MAC_0_270);
	MAC_0_271: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_271, data_out=>output_MAC_0_271);
	MAC_0_272: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_272, data_out=>output_MAC_0_272);
	MAC_0_273: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_273, data_out=>output_MAC_0_273);
	MAC_0_274: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_274, data_out=>output_MAC_0_274);
	MAC_0_275: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_275, data_out=>output_MAC_0_275);
	MAC_0_276: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_276, data_out=>output_MAC_0_276);
	MAC_0_277: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_277, data_out=>output_MAC_0_277);
	MAC_0_278: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_278, data_out=>output_MAC_0_278);
	MAC_0_279: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_279, data_out=>output_MAC_0_279);
	MAC_0_280: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_280, data_out=>output_MAC_0_280);
	MAC_0_281: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_281, data_out=>output_MAC_0_281);
	MAC_0_282: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_282, data_out=>output_MAC_0_282);
	MAC_0_283: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_283, data_out=>output_MAC_0_283);
	MAC_0_284: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_284, data_out=>output_MAC_0_284);
	MAC_0_285: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_285, data_out=>output_MAC_0_285);
	MAC_0_286: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_286, data_out=>output_MAC_0_286);
	MAC_0_287: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_287, data_out=>output_MAC_0_287);
	MAC_0_288: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_288, data_out=>output_MAC_0_288);
	MAC_0_289: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_289, data_out=>output_MAC_0_289);
	MAC_0_290: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_290, data_out=>output_MAC_0_290);
	MAC_0_291: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_291, data_out=>output_MAC_0_291);
	MAC_0_292: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_292, data_out=>output_MAC_0_292);
	MAC_0_293: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_293, data_out=>output_MAC_0_293);
	MAC_0_294: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_294, data_out=>output_MAC_0_294);
	MAC_0_295: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_295, data_out=>output_MAC_0_295);
	MAC_0_296: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_296, data_out=>output_MAC_0_296);
	MAC_0_297: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_297, data_out=>output_MAC_0_297);
	MAC_0_298: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_298, data_out=>output_MAC_0_298);
	MAC_0_299: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_299, data_out=>output_MAC_0_299);
	MAC_0_300: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_300, data_out=>output_MAC_0_300);
	MAC_0_301: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_301, data_out=>output_MAC_0_301);
	MAC_0_302: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_302, data_out=>output_MAC_0_302);
	MAC_0_303: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_303, data_out=>output_MAC_0_303);
	MAC_0_304: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_304, data_out=>output_MAC_0_304);
	MAC_0_305: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_305, data_out=>output_MAC_0_305);
	MAC_0_306: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_306, data_out=>output_MAC_0_306);
	MAC_0_307: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_307, data_out=>output_MAC_0_307);
	MAC_0_308: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_308, data_out=>output_MAC_0_308);
	MAC_0_309: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_309, data_out=>output_MAC_0_309);
	MAC_0_310: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_310, data_out=>output_MAC_0_310);
	MAC_0_311: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_311, data_out=>output_MAC_0_311);
	MAC_0_312: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_312, data_out=>output_MAC_0_312);
	MAC_0_313: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_313, data_out=>output_MAC_0_313);
	MAC_0_314: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_314, data_out=>output_MAC_0_314);
	MAC_0_315: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_315, data_out=>output_MAC_0_315);
	MAC_0_316: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_316, data_out=>output_MAC_0_316);
	MAC_0_317: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_317, data_out=>output_MAC_0_317);
	MAC_0_318: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_318, data_out=>output_MAC_0_318);
	MAC_0_319: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_319, data_out=>output_MAC_0_319);
	MAC_0_320: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_320, data_out=>output_MAC_0_320);
	MAC_0_321: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_321, data_out=>output_MAC_0_321);
	MAC_0_322: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_322, data_out=>output_MAC_0_322);
	MAC_0_323: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_323, data_out=>output_MAC_0_323);
	MAC_0_324: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_324, data_out=>output_MAC_0_324);
	MAC_0_325: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_325, data_out=>output_MAC_0_325);
	MAC_0_326: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_326, data_out=>output_MAC_0_326);
	MAC_0_327: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_327, data_out=>output_MAC_0_327);
	MAC_0_328: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_328, data_out=>output_MAC_0_328);
	MAC_0_329: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_329, data_out=>output_MAC_0_329);
	MAC_0_330: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_330, data_out=>output_MAC_0_330);
	MAC_0_331: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_331, data_out=>output_MAC_0_331);
	MAC_0_332: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_332, data_out=>output_MAC_0_332);
	MAC_0_333: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_333, data_out=>output_MAC_0_333);
	MAC_0_334: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_334, data_out=>output_MAC_0_334);
	MAC_0_335: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_335, data_out=>output_MAC_0_335);
	MAC_0_336: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_336, data_out=>output_MAC_0_336);
	MAC_0_337: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_337, data_out=>output_MAC_0_337);
	MAC_0_338: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_338, data_out=>output_MAC_0_338);
	MAC_0_339: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_339, data_out=>output_MAC_0_339);
	MAC_0_340: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_340, data_out=>output_MAC_0_340);
	MAC_0_341: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_341, data_out=>output_MAC_0_341);
	MAC_0_342: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_342, data_out=>output_MAC_0_342);
	MAC_0_343: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_343, data_out=>output_MAC_0_343);
	MAC_0_344: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_344, data_out=>output_MAC_0_344);
	MAC_0_345: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_345, data_out=>output_MAC_0_345);
	MAC_0_346: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_346, data_out=>output_MAC_0_346);
	MAC_0_347: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_347, data_out=>output_MAC_0_347);
	MAC_0_348: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_348, data_out=>output_MAC_0_348);
	MAC_0_349: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_349, data_out=>output_MAC_0_349);
	MAC_0_350: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_350, data_out=>output_MAC_0_350);
	MAC_0_351: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_351, data_out=>output_MAC_0_351);
	MAC_0_352: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_352, data_out=>output_MAC_0_352);
	MAC_0_353: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_353, data_out=>output_MAC_0_353);
	MAC_0_354: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_354, data_out=>output_MAC_0_354);
	MAC_0_355: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_355, data_out=>output_MAC_0_355);
	MAC_0_356: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_356, data_out=>output_MAC_0_356);
	MAC_0_357: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_357, data_out=>output_MAC_0_357);
	MAC_0_358: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_358, data_out=>output_MAC_0_358);
	MAC_0_359: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_359, data_out=>output_MAC_0_359);
	MAC_0_360: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_360, data_out=>output_MAC_0_360);
	MAC_0_361: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_361, data_out=>output_MAC_0_361);
	MAC_0_362: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_362, data_out=>output_MAC_0_362);
	MAC_0_363: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_363, data_out=>output_MAC_0_363);
	MAC_0_364: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_364, data_out=>output_MAC_0_364);
	MAC_0_365: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_365, data_out=>output_MAC_0_365);
	MAC_0_366: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_366, data_out=>output_MAC_0_366);
	MAC_0_367: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_367, data_out=>output_MAC_0_367);
	MAC_0_368: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_368, data_out=>output_MAC_0_368);
	MAC_0_369: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_369, data_out=>output_MAC_0_369);
	MAC_0_370: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_370, data_out=>output_MAC_0_370);
	MAC_0_371: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_371, data_out=>output_MAC_0_371);
	MAC_0_372: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_372, data_out=>output_MAC_0_372);
	MAC_0_373: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_373, data_out=>output_MAC_0_373);
	MAC_0_374: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_374, data_out=>output_MAC_0_374);
	MAC_0_375: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_375, data_out=>output_MAC_0_375);
	MAC_0_376: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_376, data_out=>output_MAC_0_376);
	MAC_0_377: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_377, data_out=>output_MAC_0_377);
	MAC_0_378: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_378, data_out=>output_MAC_0_378);
	MAC_0_379: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_379, data_out=>output_MAC_0_379);
	MAC_0_380: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_380, data_out=>output_MAC_0_380);
	MAC_0_381: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_381, data_out=>output_MAC_0_381);
	MAC_0_382: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_382, data_out=>output_MAC_0_382);
	MAC_0_383: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_383, data_out=>output_MAC_0_383);
	MAC_0_384: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_384, data_out=>output_MAC_0_384);
	MAC_0_385: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_385, data_out=>output_MAC_0_385);
	MAC_0_386: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_386, data_out=>output_MAC_0_386);
	MAC_0_387: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_387, data_out=>output_MAC_0_387);
	MAC_0_388: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_388, data_out=>output_MAC_0_388);
	MAC_0_389: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_389, data_out=>output_MAC_0_389);
	MAC_0_390: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_390, data_out=>output_MAC_0_390);
	MAC_0_391: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_391, data_out=>output_MAC_0_391);
	MAC_0_392: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_392, data_out=>output_MAC_0_392);
	MAC_0_393: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_393, data_out=>output_MAC_0_393);
	MAC_0_394: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_394, data_out=>output_MAC_0_394);
	MAC_0_395: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_395, data_out=>output_MAC_0_395);
	MAC_0_396: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_396, data_out=>output_MAC_0_396);
	MAC_0_397: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_397, data_out=>output_MAC_0_397);
	MAC_0_398: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_398, data_out=>output_MAC_0_398);
	MAC_0_399: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_399, data_out=>output_MAC_0_399);
	MAC_0_400: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_400, data_out=>output_MAC_0_400);
	MAC_0_401: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_401, data_out=>output_MAC_0_401);
	MAC_0_402: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_402, data_out=>output_MAC_0_402);
	MAC_0_403: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_403, data_out=>output_MAC_0_403);
	MAC_0_404: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_404, data_out=>output_MAC_0_404);
	MAC_0_405: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_405, data_out=>output_MAC_0_405);
	MAC_0_406: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_406, data_out=>output_MAC_0_406);
	MAC_0_407: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_407, data_out=>output_MAC_0_407);
	MAC_0_408: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_408, data_out=>output_MAC_0_408);
	MAC_0_409: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_409, data_out=>output_MAC_0_409);
	MAC_0_410: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_410, data_out=>output_MAC_0_410);
	MAC_0_411: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_411, data_out=>output_MAC_0_411);
	MAC_0_412: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_412, data_out=>output_MAC_0_412);
	MAC_0_413: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_413, data_out=>output_MAC_0_413);
	MAC_0_414: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_414, data_out=>output_MAC_0_414);
	MAC_0_415: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_415, data_out=>output_MAC_0_415);
	MAC_0_416: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_416, data_out=>output_MAC_0_416);
	MAC_0_417: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_417, data_out=>output_MAC_0_417);
	MAC_0_418: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_418, data_out=>output_MAC_0_418);
	MAC_0_419: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_419, data_out=>output_MAC_0_419);
	MAC_0_420: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_420, data_out=>output_MAC_0_420);
	MAC_0_421: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_421, data_out=>output_MAC_0_421);
	MAC_0_422: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_422, data_out=>output_MAC_0_422);
	MAC_0_423: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_423, data_out=>output_MAC_0_423);
	MAC_0_424: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_424, data_out=>output_MAC_0_424);
	MAC_0_425: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_425, data_out=>output_MAC_0_425);
	MAC_0_426: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_426, data_out=>output_MAC_0_426);
	MAC_0_427: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_427, data_out=>output_MAC_0_427);
	MAC_0_428: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_428, data_out=>output_MAC_0_428);
	MAC_0_429: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_429, data_out=>output_MAC_0_429);
	MAC_0_430: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_430, data_out=>output_MAC_0_430);
	MAC_0_431: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_431, data_out=>output_MAC_0_431);
	MAC_0_432: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_432, data_out=>output_MAC_0_432);
	MAC_0_433: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_433, data_out=>output_MAC_0_433);
	MAC_0_434: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_434, data_out=>output_MAC_0_434);
	MAC_0_435: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_435, data_out=>output_MAC_0_435);
	MAC_0_436: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_436, data_out=>output_MAC_0_436);
	MAC_0_437: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_437, data_out=>output_MAC_0_437);
	MAC_0_438: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_438, data_out=>output_MAC_0_438);
	MAC_0_439: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_439, data_out=>output_MAC_0_439);
	MAC_0_440: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_440, data_out=>output_MAC_0_440);
	MAC_0_441: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_441, data_out=>output_MAC_0_441);
	MAC_0_442: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_442, data_out=>output_MAC_0_442);
	MAC_0_443: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_443, data_out=>output_MAC_0_443);
	MAC_0_444: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_444, data_out=>output_MAC_0_444);
	MAC_0_445: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_445, data_out=>output_MAC_0_445);
	MAC_0_446: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_446, data_out=>output_MAC_0_446);
	MAC_0_447: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_447, data_out=>output_MAC_0_447);
	MAC_0_448: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_448, data_out=>output_MAC_0_448);
	MAC_0_449: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_449, data_out=>output_MAC_0_449);
	MAC_0_450: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_450, data_out=>output_MAC_0_450);
	MAC_0_451: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_451, data_out=>output_MAC_0_451);
	MAC_0_452: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_452, data_out=>output_MAC_0_452);
	MAC_0_453: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_453, data_out=>output_MAC_0_453);
	MAC_0_454: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_454, data_out=>output_MAC_0_454);
	MAC_0_455: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_455, data_out=>output_MAC_0_455);
	MAC_0_456: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_456, data_out=>output_MAC_0_456);
	MAC_0_457: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_457, data_out=>output_MAC_0_457);
	MAC_0_458: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_458, data_out=>output_MAC_0_458);
	MAC_0_459: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_459, data_out=>output_MAC_0_459);
	MAC_0_460: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_460, data_out=>output_MAC_0_460);
	MAC_0_461: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_461, data_out=>output_MAC_0_461);
	MAC_0_462: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_462, data_out=>output_MAC_0_462);
	MAC_0_463: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_463, data_out=>output_MAC_0_463);
	MAC_0_464: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_464, data_out=>output_MAC_0_464);
	MAC_0_465: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_465, data_out=>output_MAC_0_465);
	MAC_0_466: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_466, data_out=>output_MAC_0_466);
	MAC_0_467: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_467, data_out=>output_MAC_0_467);
	MAC_0_468: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_468, data_out=>output_MAC_0_468);
	MAC_0_469: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_469, data_out=>output_MAC_0_469);
	MAC_0_470: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_470, data_out=>output_MAC_0_470);
	MAC_0_471: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_471, data_out=>output_MAC_0_471);
	MAC_0_472: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_472, data_out=>output_MAC_0_472);
	MAC_0_473: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_473, data_out=>output_MAC_0_473);
	MAC_0_474: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_474, data_out=>output_MAC_0_474);
	MAC_0_475: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_475, data_out=>output_MAC_0_475);
	MAC_0_476: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_476, data_out=>output_MAC_0_476);
	MAC_0_477: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_477, data_out=>output_MAC_0_477);
	MAC_0_478: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_478, data_out=>output_MAC_0_478);
	MAC_0_479: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_479, data_out=>output_MAC_0_479);
	MAC_0_480: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_480, data_out=>output_MAC_0_480);
	MAC_0_481: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_481, data_out=>output_MAC_0_481);
	MAC_0_482: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_482, data_out=>output_MAC_0_482);
	MAC_0_483: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_483, data_out=>output_MAC_0_483);
	MAC_0_484: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_484, data_out=>output_MAC_0_484);
	MAC_0_485: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_485, data_out=>output_MAC_0_485);
	MAC_0_486: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_486, data_out=>output_MAC_0_486);
	MAC_0_487: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_487, data_out=>output_MAC_0_487);
	MAC_0_488: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_488, data_out=>output_MAC_0_488);
	MAC_0_489: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_489, data_out=>output_MAC_0_489);
	MAC_0_490: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_490, data_out=>output_MAC_0_490);
	MAC_0_491: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_491, data_out=>output_MAC_0_491);
	MAC_0_492: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_492, data_out=>output_MAC_0_492);
	MAC_0_493: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_493, data_out=>output_MAC_0_493);
	MAC_0_494: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_494, data_out=>output_MAC_0_494);
	MAC_0_495: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_495, data_out=>output_MAC_0_495);
	MAC_0_496: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_496, data_out=>output_MAC_0_496);
	MAC_0_497: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_497, data_out=>output_MAC_0_497);
	MAC_0_498: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_498, data_out=>output_MAC_0_498);
	MAC_0_499: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_499, data_out=>output_MAC_0_499);
	MAC_0_500: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_500, data_out=>output_MAC_0_500);
	MAC_0_501: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_501, data_out=>output_MAC_0_501);
	MAC_0_502: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_502, data_out=>output_MAC_0_502);
	MAC_0_503: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_503, data_out=>output_MAC_0_503);
	MAC_0_504: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_504, data_out=>output_MAC_0_504);
	MAC_0_505: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_505, data_out=>output_MAC_0_505);
	MAC_0_506: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_506, data_out=>output_MAC_0_506);
	MAC_0_507: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_507, data_out=>output_MAC_0_507);
	MAC_0_508: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_508, data_out=>output_MAC_0_508);
	MAC_0_509: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_509, data_out=>output_MAC_0_509);
	MAC_0_510: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_510, data_out=>output_MAC_0_510);
	MAC_0_511: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_511, data_out=>output_MAC_0_511);
	MAC_0_512: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_512, data_out=>output_MAC_0_512);
	MAC_0_513: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_513, data_out=>output_MAC_0_513);
	MAC_0_514: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_514, data_out=>output_MAC_0_514);
	MAC_0_515: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_515, data_out=>output_MAC_0_515);
	MAC_0_516: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_516, data_out=>output_MAC_0_516);
	MAC_0_517: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_517, data_out=>output_MAC_0_517);
	MAC_0_518: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_518, data_out=>output_MAC_0_518);
	MAC_0_519: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_519, data_out=>output_MAC_0_519);
	MAC_0_520: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_520, data_out=>output_MAC_0_520);
	MAC_0_521: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_521, data_out=>output_MAC_0_521);
	MAC_0_522: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_522, data_out=>output_MAC_0_522);
	MAC_0_523: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_523, data_out=>output_MAC_0_523);
	MAC_0_524: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_524, data_out=>output_MAC_0_524);
	MAC_0_525: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_525, data_out=>output_MAC_0_525);
	MAC_0_526: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_526, data_out=>output_MAC_0_526);
	MAC_0_527: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_527, data_out=>output_MAC_0_527);
	MAC_0_528: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_528, data_out=>output_MAC_0_528);
	MAC_0_529: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_529, data_out=>output_MAC_0_529);
	MAC_0_530: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_530, data_out=>output_MAC_0_530);
	MAC_0_531: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_531, data_out=>output_MAC_0_531);
	MAC_0_532: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_532, data_out=>output_MAC_0_532);
	MAC_0_533: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_533, data_out=>output_MAC_0_533);
	MAC_0_534: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_534, data_out=>output_MAC_0_534);
	MAC_0_535: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_535, data_out=>output_MAC_0_535);
	MAC_0_536: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_536, data_out=>output_MAC_0_536);
	MAC_0_537: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_537, data_out=>output_MAC_0_537);
	MAC_0_538: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_538, data_out=>output_MAC_0_538);
	MAC_0_539: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_539, data_out=>output_MAC_0_539);
	MAC_0_540: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_540, data_out=>output_MAC_0_540);
	MAC_0_541: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_541, data_out=>output_MAC_0_541);
	MAC_0_542: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_542, data_out=>output_MAC_0_542);
	MAC_0_543: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_543, data_out=>output_MAC_0_543);
	MAC_0_544: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_544, data_out=>output_MAC_0_544);
	MAC_0_545: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_545, data_out=>output_MAC_0_545);
	MAC_0_546: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_546, data_out=>output_MAC_0_546);
	MAC_0_547: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_547, data_out=>output_MAC_0_547);
	MAC_0_548: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_548, data_out=>output_MAC_0_548);
	MAC_0_549: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_549, data_out=>output_MAC_0_549);
	MAC_0_550: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_550, data_out=>output_MAC_0_550);
	MAC_0_551: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_551, data_out=>output_MAC_0_551);
	MAC_0_552: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_552, data_out=>output_MAC_0_552);
	MAC_0_553: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_553, data_out=>output_MAC_0_553);
	MAC_0_554: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_554, data_out=>output_MAC_0_554);
	MAC_0_555: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_555, data_out=>output_MAC_0_555);
	MAC_0_556: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_556, data_out=>output_MAC_0_556);
	MAC_0_557: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_557, data_out=>output_MAC_0_557);
	MAC_0_558: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_558, data_out=>output_MAC_0_558);
	MAC_0_559: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_559, data_out=>output_MAC_0_559);
	MAC_0_560: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_560, data_out=>output_MAC_0_560);
	MAC_0_561: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_561, data_out=>output_MAC_0_561);
	MAC_0_562: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_562, data_out=>output_MAC_0_562);
	MAC_0_563: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_563, data_out=>output_MAC_0_563);
	MAC_0_564: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_564, data_out=>output_MAC_0_564);
	MAC_0_565: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_565, data_out=>output_MAC_0_565);
	MAC_0_566: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_566, data_out=>output_MAC_0_566);
	MAC_0_567: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_567, data_out=>output_MAC_0_567);
	MAC_0_568: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_568, data_out=>output_MAC_0_568);
	MAC_0_569: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_569, data_out=>output_MAC_0_569);
	MAC_0_570: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_570, data_out=>output_MAC_0_570);
	MAC_0_571: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_571, data_out=>output_MAC_0_571);
	MAC_0_572: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_572, data_out=>output_MAC_0_572);
	MAC_0_573: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_573, data_out=>output_MAC_0_573);
	MAC_0_574: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_574, data_out=>output_MAC_0_574);
	MAC_0_575: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_575, data_out=>output_MAC_0_575);
	MAC_0_576: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_576, data_out=>output_MAC_0_576);
	MAC_0_577: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_577, data_out=>output_MAC_0_577);
	MAC_0_578: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_578, data_out=>output_MAC_0_578);
	MAC_0_579: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_579, data_out=>output_MAC_0_579);
	MAC_0_580: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_580, data_out=>output_MAC_0_580);
	MAC_0_581: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_581, data_out=>output_MAC_0_581);
	MAC_0_582: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_582, data_out=>output_MAC_0_582);
	MAC_0_583: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_583, data_out=>output_MAC_0_583);
	MAC_0_584: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_584, data_out=>output_MAC_0_584);
	MAC_0_585: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_585, data_out=>output_MAC_0_585);
	MAC_0_586: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_586, data_out=>output_MAC_0_586);
	MAC_0_587: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_587, data_out=>output_MAC_0_587);
	MAC_0_588: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_588, data_out=>output_MAC_0_588);
	MAC_0_589: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_589, data_out=>output_MAC_0_589);
	MAC_0_590: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_590, data_out=>output_MAC_0_590);
	MAC_0_591: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_591, data_out=>output_MAC_0_591);
	MAC_0_592: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_592, data_out=>output_MAC_0_592);
	MAC_0_593: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_593, data_out=>output_MAC_0_593);
	MAC_0_594: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_594, data_out=>output_MAC_0_594);
	MAC_0_595: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_595, data_out=>output_MAC_0_595);
	MAC_0_596: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_596, data_out=>output_MAC_0_596);
	MAC_0_597: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_597, data_out=>output_MAC_0_597);
	MAC_0_598: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_598, data_out=>output_MAC_0_598);
	MAC_0_599: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_599, data_out=>output_MAC_0_599);
	MAC_0_600: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_600, data_out=>output_MAC_0_600);
	MAC_0_601: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_601, data_out=>output_MAC_0_601);
	MAC_0_602: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_602, data_out=>output_MAC_0_602);
	MAC_0_603: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_603, data_out=>output_MAC_0_603);
	MAC_0_604: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_604, data_out=>output_MAC_0_604);
	MAC_0_605: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_605, data_out=>output_MAC_0_605);
	MAC_0_606: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_606, data_out=>output_MAC_0_606);
	MAC_0_607: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_607, data_out=>output_MAC_0_607);
	MAC_0_608: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_608, data_out=>output_MAC_0_608);
	MAC_0_609: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_609, data_out=>output_MAC_0_609);
	MAC_0_610: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_610, data_out=>output_MAC_0_610);
	MAC_0_611: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_611, data_out=>output_MAC_0_611);
	MAC_0_612: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_612, data_out=>output_MAC_0_612);
	MAC_0_613: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_613, data_out=>output_MAC_0_613);
	MAC_0_614: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_614, data_out=>output_MAC_0_614);
	MAC_0_615: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_615, data_out=>output_MAC_0_615);
	MAC_0_616: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_616, data_out=>output_MAC_0_616);
	MAC_0_617: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_617, data_out=>output_MAC_0_617);
	MAC_0_618: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_618, data_out=>output_MAC_0_618);
	MAC_0_619: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_619, data_out=>output_MAC_0_619);
	MAC_0_620: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_620, data_out=>output_MAC_0_620);
	MAC_0_621: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_621, data_out=>output_MAC_0_621);
	MAC_0_622: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_622, data_out=>output_MAC_0_622);
	MAC_0_623: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_623, data_out=>output_MAC_0_623);
	MAC_0_624: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_624, data_out=>output_MAC_0_624);
	MAC_0_625: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_625, data_out=>output_MAC_0_625);
	MAC_0_626: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_626, data_out=>output_MAC_0_626);
	MAC_0_627: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_627, data_out=>output_MAC_0_627);
	MAC_0_628: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_628, data_out=>output_MAC_0_628);
	MAC_0_629: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_629, data_out=>output_MAC_0_629);
	MAC_0_630: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_630, data_out=>output_MAC_0_630);
	MAC_0_631: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_631, data_out=>output_MAC_0_631);
	MAC_0_632: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_632, data_out=>output_MAC_0_632);
	MAC_0_633: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_633, data_out=>output_MAC_0_633);
	MAC_0_634: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_634, data_out=>output_MAC_0_634);
	MAC_0_635: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_635, data_out=>output_MAC_0_635);
	MAC_0_636: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_636, data_out=>output_MAC_0_636);
	MAC_0_637: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_637, data_out=>output_MAC_0_637);
	MAC_0_638: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_638, data_out=>output_MAC_0_638);
	MAC_0_639: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_639, data_out=>output_MAC_0_639);
	MAC_0_640: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_640, data_out=>output_MAC_0_640);
	MAC_0_641: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_641, data_out=>output_MAC_0_641);
	MAC_0_642: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_642, data_out=>output_MAC_0_642);
	MAC_0_643: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_643, data_out=>output_MAC_0_643);
	MAC_0_644: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_644, data_out=>output_MAC_0_644);
	MAC_0_645: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_645, data_out=>output_MAC_0_645);
	MAC_0_646: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_646, data_out=>output_MAC_0_646);
	MAC_0_647: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_647, data_out=>output_MAC_0_647);
	MAC_0_648: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_648, data_out=>output_MAC_0_648);
	MAC_0_649: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_649, data_out=>output_MAC_0_649);
	MAC_0_650: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_650, data_out=>output_MAC_0_650);
	MAC_0_651: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_651, data_out=>output_MAC_0_651);
	MAC_0_652: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_652, data_out=>output_MAC_0_652);
	MAC_0_653: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_653, data_out=>output_MAC_0_653);
	MAC_0_654: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_654, data_out=>output_MAC_0_654);
	MAC_0_655: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_655, data_out=>output_MAC_0_655);
	MAC_0_656: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_656, data_out=>output_MAC_0_656);
	MAC_0_657: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_657, data_out=>output_MAC_0_657);
	MAC_0_658: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_658, data_out=>output_MAC_0_658);
	MAC_0_659: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_659, data_out=>output_MAC_0_659);
	MAC_0_660: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_660, data_out=>output_MAC_0_660);
	MAC_0_661: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_661, data_out=>output_MAC_0_661);
	MAC_0_662: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_662, data_out=>output_MAC_0_662);
	MAC_0_663: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_663, data_out=>output_MAC_0_663);
	MAC_0_664: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_664, data_out=>output_MAC_0_664);
	MAC_0_665: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_665, data_out=>output_MAC_0_665);
	MAC_0_666: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_666, data_out=>output_MAC_0_666);
	MAC_0_667: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_667, data_out=>output_MAC_0_667);
	MAC_0_668: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_668, data_out=>output_MAC_0_668);
	MAC_0_669: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_669, data_out=>output_MAC_0_669);
	MAC_0_670: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_670, data_out=>output_MAC_0_670);
	MAC_0_671: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_671, data_out=>output_MAC_0_671);
	MAC_0_672: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_672, data_out=>output_MAC_0_672);
	MAC_0_673: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_673, data_out=>output_MAC_0_673);
	MAC_0_674: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_674, data_out=>output_MAC_0_674);
	MAC_0_675: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_675, data_out=>output_MAC_0_675);
	MAC_0_676: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_676, data_out=>output_MAC_0_676);
	MAC_0_677: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_677, data_out=>output_MAC_0_677);
	MAC_0_678: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_678, data_out=>output_MAC_0_678);
	MAC_0_679: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_679, data_out=>output_MAC_0_679);
	MAC_0_680: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_680, data_out=>output_MAC_0_680);
	MAC_0_681: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_681, data_out=>output_MAC_0_681);
	MAC_0_682: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_682, data_out=>output_MAC_0_682);
	MAC_0_683: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_683, data_out=>output_MAC_0_683);
	MAC_0_684: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_684, data_out=>output_MAC_0_684);
	MAC_0_685: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_685, data_out=>output_MAC_0_685);
	MAC_0_686: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_686, data_out=>output_MAC_0_686);
	MAC_0_687: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_687, data_out=>output_MAC_0_687);
	MAC_0_688: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_688, data_out=>output_MAC_0_688);
	MAC_0_689: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_689, data_out=>output_MAC_0_689);
	MAC_0_690: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_690, data_out=>output_MAC_0_690);
	MAC_0_691: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_691, data_out=>output_MAC_0_691);
	MAC_0_692: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_692, data_out=>output_MAC_0_692);
	MAC_0_693: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_693, data_out=>output_MAC_0_693);
	MAC_0_694: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_694, data_out=>output_MAC_0_694);
	MAC_0_695: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_695, data_out=>output_MAC_0_695);
	MAC_0_696: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_696, data_out=>output_MAC_0_696);
	MAC_0_697: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_697, data_out=>output_MAC_0_697);
	MAC_0_698: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_698, data_out=>output_MAC_0_698);
	MAC_0_699: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_699, data_out=>output_MAC_0_699);
	MAC_0_700: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_700, data_out=>output_MAC_0_700);
	MAC_0_701: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_701, data_out=>output_MAC_0_701);
	MAC_0_702: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_702, data_out=>output_MAC_0_702);
	MAC_0_703: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_703, data_out=>output_MAC_0_703);
	MAC_0_704: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_704, data_out=>output_MAC_0_704);
	MAC_0_705: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_705, data_out=>output_MAC_0_705);
	MAC_0_706: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_706, data_out=>output_MAC_0_706);
	MAC_0_707: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_707, data_out=>output_MAC_0_707);
	MAC_0_708: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_708, data_out=>output_MAC_0_708);
	MAC_0_709: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_709, data_out=>output_MAC_0_709);
	MAC_0_710: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_710, data_out=>output_MAC_0_710);
	MAC_0_711: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_711, data_out=>output_MAC_0_711);
	MAC_0_712: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_712, data_out=>output_MAC_0_712);
	MAC_0_713: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_713, data_out=>output_MAC_0_713);
	MAC_0_714: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_714, data_out=>output_MAC_0_714);
	MAC_0_715: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_715, data_out=>output_MAC_0_715);
	MAC_0_716: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_716, data_out=>output_MAC_0_716);
	MAC_0_717: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_717, data_out=>output_MAC_0_717);
	MAC_0_718: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_718, data_out=>output_MAC_0_718);
	MAC_0_719: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_719, data_out=>output_MAC_0_719);
	MAC_0_720: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_720, data_out=>output_MAC_0_720);
	MAC_0_721: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_721, data_out=>output_MAC_0_721);
	MAC_0_722: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_722, data_out=>output_MAC_0_722);
	MAC_0_723: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_723, data_out=>output_MAC_0_723);
	MAC_0_724: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_724, data_out=>output_MAC_0_724);
	MAC_0_725: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_725, data_out=>output_MAC_0_725);
	MAC_0_726: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_726, data_out=>output_MAC_0_726);
	MAC_0_727: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_727, data_out=>output_MAC_0_727);
	MAC_0_728: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_728, data_out=>output_MAC_0_728);
	MAC_0_729: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_729, data_out=>output_MAC_0_729);
	MAC_0_730: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_730, data_out=>output_MAC_0_730);
	MAC_0_731: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_731, data_out=>output_MAC_0_731);
	MAC_0_732: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_732, data_out=>output_MAC_0_732);
	MAC_0_733: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_733, data_out=>output_MAC_0_733);
	MAC_0_734: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_734, data_out=>output_MAC_0_734);
	MAC_0_735: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_735, data_out=>output_MAC_0_735);
	MAC_0_736: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_736, data_out=>output_MAC_0_736);
	MAC_0_737: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_737, data_out=>output_MAC_0_737);
	MAC_0_738: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_738, data_out=>output_MAC_0_738);
	MAC_0_739: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_739, data_out=>output_MAC_0_739);
	MAC_0_740: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_740, data_out=>output_MAC_0_740);
	MAC_0_741: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_741, data_out=>output_MAC_0_741);
	MAC_0_742: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_742, data_out=>output_MAC_0_742);
	MAC_0_743: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_743, data_out=>output_MAC_0_743);
	MAC_0_744: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_744, data_out=>output_MAC_0_744);
	MAC_0_745: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_745, data_out=>output_MAC_0_745);
	MAC_0_746: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_746, data_out=>output_MAC_0_746);
	MAC_0_747: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_747, data_out=>output_MAC_0_747);
	MAC_0_748: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_748, data_out=>output_MAC_0_748);
	MAC_0_749: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_749, data_out=>output_MAC_0_749);
	MAC_0_750: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_750, data_out=>output_MAC_0_750);
	MAC_0_751: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_751, data_out=>output_MAC_0_751);
	MAC_0_752: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_752, data_out=>output_MAC_0_752);
	MAC_0_753: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_753, data_out=>output_MAC_0_753);
	MAC_0_754: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_754, data_out=>output_MAC_0_754);
	MAC_0_755: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_755, data_out=>output_MAC_0_755);
	MAC_0_756: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_756, data_out=>output_MAC_0_756);
	MAC_0_757: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_757, data_out=>output_MAC_0_757);
	MAC_0_758: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_758, data_out=>output_MAC_0_758);
	MAC_0_759: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_759, data_out=>output_MAC_0_759);
	MAC_0_760: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_760, data_out=>output_MAC_0_760);
	MAC_0_761: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_761, data_out=>output_MAC_0_761);
	MAC_0_762: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_762, data_out=>output_MAC_0_762);
	MAC_0_763: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_763, data_out=>output_MAC_0_763);
	MAC_0_764: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_764, data_out=>output_MAC_0_764);
	MAC_0_765: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_765, data_out=>output_MAC_0_765);
	MAC_0_766: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_766, data_out=>output_MAC_0_766);
	MAC_0_767: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_0, data_in_B=>input_col_767, data_out=>output_MAC_0_767);
	MAC_1_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_0, data_out=>output_MAC_1_0);
	MAC_1_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_1, data_out=>output_MAC_1_1);
	MAC_1_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_2, data_out=>output_MAC_1_2);
	MAC_1_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_3, data_out=>output_MAC_1_3);
	MAC_1_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_4, data_out=>output_MAC_1_4);
	MAC_1_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_5, data_out=>output_MAC_1_5);
	MAC_1_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_6, data_out=>output_MAC_1_6);
	MAC_1_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_7, data_out=>output_MAC_1_7);
	MAC_1_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_8, data_out=>output_MAC_1_8);
	MAC_1_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_9, data_out=>output_MAC_1_9);
	MAC_1_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_10, data_out=>output_MAC_1_10);
	MAC_1_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_11, data_out=>output_MAC_1_11);
	MAC_1_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_12, data_out=>output_MAC_1_12);
	MAC_1_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_13, data_out=>output_MAC_1_13);
	MAC_1_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_14, data_out=>output_MAC_1_14);
	MAC_1_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_15, data_out=>output_MAC_1_15);
	MAC_1_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_16, data_out=>output_MAC_1_16);
	MAC_1_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_17, data_out=>output_MAC_1_17);
	MAC_1_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_18, data_out=>output_MAC_1_18);
	MAC_1_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_19, data_out=>output_MAC_1_19);
	MAC_1_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_20, data_out=>output_MAC_1_20);
	MAC_1_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_21, data_out=>output_MAC_1_21);
	MAC_1_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_22, data_out=>output_MAC_1_22);
	MAC_1_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_23, data_out=>output_MAC_1_23);
	MAC_1_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_24, data_out=>output_MAC_1_24);
	MAC_1_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_25, data_out=>output_MAC_1_25);
	MAC_1_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_26, data_out=>output_MAC_1_26);
	MAC_1_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_27, data_out=>output_MAC_1_27);
	MAC_1_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_28, data_out=>output_MAC_1_28);
	MAC_1_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_29, data_out=>output_MAC_1_29);
	MAC_1_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_30, data_out=>output_MAC_1_30);
	MAC_1_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_31, data_out=>output_MAC_1_31);
	MAC_1_32: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_32, data_out=>output_MAC_1_32);
	MAC_1_33: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_33, data_out=>output_MAC_1_33);
	MAC_1_34: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_34, data_out=>output_MAC_1_34);
	MAC_1_35: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_35, data_out=>output_MAC_1_35);
	MAC_1_36: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_36, data_out=>output_MAC_1_36);
	MAC_1_37: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_37, data_out=>output_MAC_1_37);
	MAC_1_38: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_38, data_out=>output_MAC_1_38);
	MAC_1_39: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_39, data_out=>output_MAC_1_39);
	MAC_1_40: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_40, data_out=>output_MAC_1_40);
	MAC_1_41: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_41, data_out=>output_MAC_1_41);
	MAC_1_42: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_42, data_out=>output_MAC_1_42);
	MAC_1_43: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_43, data_out=>output_MAC_1_43);
	MAC_1_44: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_44, data_out=>output_MAC_1_44);
	MAC_1_45: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_45, data_out=>output_MAC_1_45);
	MAC_1_46: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_46, data_out=>output_MAC_1_46);
	MAC_1_47: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_47, data_out=>output_MAC_1_47);
	MAC_1_48: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_48, data_out=>output_MAC_1_48);
	MAC_1_49: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_49, data_out=>output_MAC_1_49);
	MAC_1_50: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_50, data_out=>output_MAC_1_50);
	MAC_1_51: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_51, data_out=>output_MAC_1_51);
	MAC_1_52: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_52, data_out=>output_MAC_1_52);
	MAC_1_53: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_53, data_out=>output_MAC_1_53);
	MAC_1_54: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_54, data_out=>output_MAC_1_54);
	MAC_1_55: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_55, data_out=>output_MAC_1_55);
	MAC_1_56: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_56, data_out=>output_MAC_1_56);
	MAC_1_57: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_57, data_out=>output_MAC_1_57);
	MAC_1_58: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_58, data_out=>output_MAC_1_58);
	MAC_1_59: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_59, data_out=>output_MAC_1_59);
	MAC_1_60: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_60, data_out=>output_MAC_1_60);
	MAC_1_61: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_61, data_out=>output_MAC_1_61);
	MAC_1_62: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_62, data_out=>output_MAC_1_62);
	MAC_1_63: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_63, data_out=>output_MAC_1_63);
	MAC_1_64: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_64, data_out=>output_MAC_1_64);
	MAC_1_65: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_65, data_out=>output_MAC_1_65);
	MAC_1_66: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_66, data_out=>output_MAC_1_66);
	MAC_1_67: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_67, data_out=>output_MAC_1_67);
	MAC_1_68: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_68, data_out=>output_MAC_1_68);
	MAC_1_69: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_69, data_out=>output_MAC_1_69);
	MAC_1_70: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_70, data_out=>output_MAC_1_70);
	MAC_1_71: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_71, data_out=>output_MAC_1_71);
	MAC_1_72: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_72, data_out=>output_MAC_1_72);
	MAC_1_73: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_73, data_out=>output_MAC_1_73);
	MAC_1_74: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_74, data_out=>output_MAC_1_74);
	MAC_1_75: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_75, data_out=>output_MAC_1_75);
	MAC_1_76: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_76, data_out=>output_MAC_1_76);
	MAC_1_77: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_77, data_out=>output_MAC_1_77);
	MAC_1_78: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_78, data_out=>output_MAC_1_78);
	MAC_1_79: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_79, data_out=>output_MAC_1_79);
	MAC_1_80: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_80, data_out=>output_MAC_1_80);
	MAC_1_81: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_81, data_out=>output_MAC_1_81);
	MAC_1_82: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_82, data_out=>output_MAC_1_82);
	MAC_1_83: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_83, data_out=>output_MAC_1_83);
	MAC_1_84: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_84, data_out=>output_MAC_1_84);
	MAC_1_85: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_85, data_out=>output_MAC_1_85);
	MAC_1_86: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_86, data_out=>output_MAC_1_86);
	MAC_1_87: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_87, data_out=>output_MAC_1_87);
	MAC_1_88: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_88, data_out=>output_MAC_1_88);
	MAC_1_89: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_89, data_out=>output_MAC_1_89);
	MAC_1_90: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_90, data_out=>output_MAC_1_90);
	MAC_1_91: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_91, data_out=>output_MAC_1_91);
	MAC_1_92: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_92, data_out=>output_MAC_1_92);
	MAC_1_93: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_93, data_out=>output_MAC_1_93);
	MAC_1_94: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_94, data_out=>output_MAC_1_94);
	MAC_1_95: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_95, data_out=>output_MAC_1_95);
	MAC_1_96: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_96, data_out=>output_MAC_1_96);
	MAC_1_97: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_97, data_out=>output_MAC_1_97);
	MAC_1_98: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_98, data_out=>output_MAC_1_98);
	MAC_1_99: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_99, data_out=>output_MAC_1_99);
	MAC_1_100: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_100, data_out=>output_MAC_1_100);
	MAC_1_101: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_101, data_out=>output_MAC_1_101);
	MAC_1_102: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_102, data_out=>output_MAC_1_102);
	MAC_1_103: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_103, data_out=>output_MAC_1_103);
	MAC_1_104: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_104, data_out=>output_MAC_1_104);
	MAC_1_105: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_105, data_out=>output_MAC_1_105);
	MAC_1_106: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_106, data_out=>output_MAC_1_106);
	MAC_1_107: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_107, data_out=>output_MAC_1_107);
	MAC_1_108: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_108, data_out=>output_MAC_1_108);
	MAC_1_109: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_109, data_out=>output_MAC_1_109);
	MAC_1_110: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_110, data_out=>output_MAC_1_110);
	MAC_1_111: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_111, data_out=>output_MAC_1_111);
	MAC_1_112: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_112, data_out=>output_MAC_1_112);
	MAC_1_113: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_113, data_out=>output_MAC_1_113);
	MAC_1_114: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_114, data_out=>output_MAC_1_114);
	MAC_1_115: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_115, data_out=>output_MAC_1_115);
	MAC_1_116: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_116, data_out=>output_MAC_1_116);
	MAC_1_117: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_117, data_out=>output_MAC_1_117);
	MAC_1_118: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_118, data_out=>output_MAC_1_118);
	MAC_1_119: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_119, data_out=>output_MAC_1_119);
	MAC_1_120: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_120, data_out=>output_MAC_1_120);
	MAC_1_121: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_121, data_out=>output_MAC_1_121);
	MAC_1_122: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_122, data_out=>output_MAC_1_122);
	MAC_1_123: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_123, data_out=>output_MAC_1_123);
	MAC_1_124: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_124, data_out=>output_MAC_1_124);
	MAC_1_125: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_125, data_out=>output_MAC_1_125);
	MAC_1_126: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_126, data_out=>output_MAC_1_126);
	MAC_1_127: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_127, data_out=>output_MAC_1_127);
	MAC_1_128: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_128, data_out=>output_MAC_1_128);
	MAC_1_129: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_129, data_out=>output_MAC_1_129);
	MAC_1_130: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_130, data_out=>output_MAC_1_130);
	MAC_1_131: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_131, data_out=>output_MAC_1_131);
	MAC_1_132: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_132, data_out=>output_MAC_1_132);
	MAC_1_133: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_133, data_out=>output_MAC_1_133);
	MAC_1_134: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_134, data_out=>output_MAC_1_134);
	MAC_1_135: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_135, data_out=>output_MAC_1_135);
	MAC_1_136: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_136, data_out=>output_MAC_1_136);
	MAC_1_137: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_137, data_out=>output_MAC_1_137);
	MAC_1_138: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_138, data_out=>output_MAC_1_138);
	MAC_1_139: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_139, data_out=>output_MAC_1_139);
	MAC_1_140: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_140, data_out=>output_MAC_1_140);
	MAC_1_141: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_141, data_out=>output_MAC_1_141);
	MAC_1_142: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_142, data_out=>output_MAC_1_142);
	MAC_1_143: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_143, data_out=>output_MAC_1_143);
	MAC_1_144: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_144, data_out=>output_MAC_1_144);
	MAC_1_145: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_145, data_out=>output_MAC_1_145);
	MAC_1_146: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_146, data_out=>output_MAC_1_146);
	MAC_1_147: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_147, data_out=>output_MAC_1_147);
	MAC_1_148: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_148, data_out=>output_MAC_1_148);
	MAC_1_149: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_149, data_out=>output_MAC_1_149);
	MAC_1_150: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_150, data_out=>output_MAC_1_150);
	MAC_1_151: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_151, data_out=>output_MAC_1_151);
	MAC_1_152: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_152, data_out=>output_MAC_1_152);
	MAC_1_153: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_153, data_out=>output_MAC_1_153);
	MAC_1_154: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_154, data_out=>output_MAC_1_154);
	MAC_1_155: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_155, data_out=>output_MAC_1_155);
	MAC_1_156: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_156, data_out=>output_MAC_1_156);
	MAC_1_157: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_157, data_out=>output_MAC_1_157);
	MAC_1_158: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_158, data_out=>output_MAC_1_158);
	MAC_1_159: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_159, data_out=>output_MAC_1_159);
	MAC_1_160: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_160, data_out=>output_MAC_1_160);
	MAC_1_161: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_161, data_out=>output_MAC_1_161);
	MAC_1_162: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_162, data_out=>output_MAC_1_162);
	MAC_1_163: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_163, data_out=>output_MAC_1_163);
	MAC_1_164: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_164, data_out=>output_MAC_1_164);
	MAC_1_165: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_165, data_out=>output_MAC_1_165);
	MAC_1_166: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_166, data_out=>output_MAC_1_166);
	MAC_1_167: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_167, data_out=>output_MAC_1_167);
	MAC_1_168: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_168, data_out=>output_MAC_1_168);
	MAC_1_169: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_169, data_out=>output_MAC_1_169);
	MAC_1_170: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_170, data_out=>output_MAC_1_170);
	MAC_1_171: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_171, data_out=>output_MAC_1_171);
	MAC_1_172: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_172, data_out=>output_MAC_1_172);
	MAC_1_173: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_173, data_out=>output_MAC_1_173);
	MAC_1_174: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_174, data_out=>output_MAC_1_174);
	MAC_1_175: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_175, data_out=>output_MAC_1_175);
	MAC_1_176: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_176, data_out=>output_MAC_1_176);
	MAC_1_177: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_177, data_out=>output_MAC_1_177);
	MAC_1_178: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_178, data_out=>output_MAC_1_178);
	MAC_1_179: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_179, data_out=>output_MAC_1_179);
	MAC_1_180: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_180, data_out=>output_MAC_1_180);
	MAC_1_181: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_181, data_out=>output_MAC_1_181);
	MAC_1_182: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_182, data_out=>output_MAC_1_182);
	MAC_1_183: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_183, data_out=>output_MAC_1_183);
	MAC_1_184: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_184, data_out=>output_MAC_1_184);
	MAC_1_185: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_185, data_out=>output_MAC_1_185);
	MAC_1_186: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_186, data_out=>output_MAC_1_186);
	MAC_1_187: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_187, data_out=>output_MAC_1_187);
	MAC_1_188: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_188, data_out=>output_MAC_1_188);
	MAC_1_189: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_189, data_out=>output_MAC_1_189);
	MAC_1_190: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_190, data_out=>output_MAC_1_190);
	MAC_1_191: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_191, data_out=>output_MAC_1_191);
	MAC_1_192: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_192, data_out=>output_MAC_1_192);
	MAC_1_193: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_193, data_out=>output_MAC_1_193);
	MAC_1_194: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_194, data_out=>output_MAC_1_194);
	MAC_1_195: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_195, data_out=>output_MAC_1_195);
	MAC_1_196: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_196, data_out=>output_MAC_1_196);
	MAC_1_197: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_197, data_out=>output_MAC_1_197);
	MAC_1_198: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_198, data_out=>output_MAC_1_198);
	MAC_1_199: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_199, data_out=>output_MAC_1_199);
	MAC_1_200: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_200, data_out=>output_MAC_1_200);
	MAC_1_201: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_201, data_out=>output_MAC_1_201);
	MAC_1_202: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_202, data_out=>output_MAC_1_202);
	MAC_1_203: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_203, data_out=>output_MAC_1_203);
	MAC_1_204: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_204, data_out=>output_MAC_1_204);
	MAC_1_205: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_205, data_out=>output_MAC_1_205);
	MAC_1_206: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_206, data_out=>output_MAC_1_206);
	MAC_1_207: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_207, data_out=>output_MAC_1_207);
	MAC_1_208: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_208, data_out=>output_MAC_1_208);
	MAC_1_209: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_209, data_out=>output_MAC_1_209);
	MAC_1_210: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_210, data_out=>output_MAC_1_210);
	MAC_1_211: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_211, data_out=>output_MAC_1_211);
	MAC_1_212: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_212, data_out=>output_MAC_1_212);
	MAC_1_213: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_213, data_out=>output_MAC_1_213);
	MAC_1_214: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_214, data_out=>output_MAC_1_214);
	MAC_1_215: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_215, data_out=>output_MAC_1_215);
	MAC_1_216: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_216, data_out=>output_MAC_1_216);
	MAC_1_217: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_217, data_out=>output_MAC_1_217);
	MAC_1_218: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_218, data_out=>output_MAC_1_218);
	MAC_1_219: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_219, data_out=>output_MAC_1_219);
	MAC_1_220: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_220, data_out=>output_MAC_1_220);
	MAC_1_221: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_221, data_out=>output_MAC_1_221);
	MAC_1_222: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_222, data_out=>output_MAC_1_222);
	MAC_1_223: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_223, data_out=>output_MAC_1_223);
	MAC_1_224: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_224, data_out=>output_MAC_1_224);
	MAC_1_225: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_225, data_out=>output_MAC_1_225);
	MAC_1_226: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_226, data_out=>output_MAC_1_226);
	MAC_1_227: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_227, data_out=>output_MAC_1_227);
	MAC_1_228: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_228, data_out=>output_MAC_1_228);
	MAC_1_229: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_229, data_out=>output_MAC_1_229);
	MAC_1_230: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_230, data_out=>output_MAC_1_230);
	MAC_1_231: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_231, data_out=>output_MAC_1_231);
	MAC_1_232: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_232, data_out=>output_MAC_1_232);
	MAC_1_233: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_233, data_out=>output_MAC_1_233);
	MAC_1_234: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_234, data_out=>output_MAC_1_234);
	MAC_1_235: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_235, data_out=>output_MAC_1_235);
	MAC_1_236: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_236, data_out=>output_MAC_1_236);
	MAC_1_237: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_237, data_out=>output_MAC_1_237);
	MAC_1_238: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_238, data_out=>output_MAC_1_238);
	MAC_1_239: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_239, data_out=>output_MAC_1_239);
	MAC_1_240: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_240, data_out=>output_MAC_1_240);
	MAC_1_241: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_241, data_out=>output_MAC_1_241);
	MAC_1_242: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_242, data_out=>output_MAC_1_242);
	MAC_1_243: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_243, data_out=>output_MAC_1_243);
	MAC_1_244: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_244, data_out=>output_MAC_1_244);
	MAC_1_245: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_245, data_out=>output_MAC_1_245);
	MAC_1_246: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_246, data_out=>output_MAC_1_246);
	MAC_1_247: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_247, data_out=>output_MAC_1_247);
	MAC_1_248: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_248, data_out=>output_MAC_1_248);
	MAC_1_249: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_249, data_out=>output_MAC_1_249);
	MAC_1_250: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_250, data_out=>output_MAC_1_250);
	MAC_1_251: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_251, data_out=>output_MAC_1_251);
	MAC_1_252: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_252, data_out=>output_MAC_1_252);
	MAC_1_253: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_253, data_out=>output_MAC_1_253);
	MAC_1_254: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_254, data_out=>output_MAC_1_254);
	MAC_1_255: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_255, data_out=>output_MAC_1_255);
	MAC_1_256: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_256, data_out=>output_MAC_1_256);
	MAC_1_257: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_257, data_out=>output_MAC_1_257);
	MAC_1_258: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_258, data_out=>output_MAC_1_258);
	MAC_1_259: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_259, data_out=>output_MAC_1_259);
	MAC_1_260: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_260, data_out=>output_MAC_1_260);
	MAC_1_261: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_261, data_out=>output_MAC_1_261);
	MAC_1_262: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_262, data_out=>output_MAC_1_262);
	MAC_1_263: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_263, data_out=>output_MAC_1_263);
	MAC_1_264: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_264, data_out=>output_MAC_1_264);
	MAC_1_265: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_265, data_out=>output_MAC_1_265);
	MAC_1_266: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_266, data_out=>output_MAC_1_266);
	MAC_1_267: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_267, data_out=>output_MAC_1_267);
	MAC_1_268: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_268, data_out=>output_MAC_1_268);
	MAC_1_269: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_269, data_out=>output_MAC_1_269);
	MAC_1_270: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_270, data_out=>output_MAC_1_270);
	MAC_1_271: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_271, data_out=>output_MAC_1_271);
	MAC_1_272: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_272, data_out=>output_MAC_1_272);
	MAC_1_273: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_273, data_out=>output_MAC_1_273);
	MAC_1_274: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_274, data_out=>output_MAC_1_274);
	MAC_1_275: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_275, data_out=>output_MAC_1_275);
	MAC_1_276: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_276, data_out=>output_MAC_1_276);
	MAC_1_277: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_277, data_out=>output_MAC_1_277);
	MAC_1_278: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_278, data_out=>output_MAC_1_278);
	MAC_1_279: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_279, data_out=>output_MAC_1_279);
	MAC_1_280: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_280, data_out=>output_MAC_1_280);
	MAC_1_281: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_281, data_out=>output_MAC_1_281);
	MAC_1_282: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_282, data_out=>output_MAC_1_282);
	MAC_1_283: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_283, data_out=>output_MAC_1_283);
	MAC_1_284: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_284, data_out=>output_MAC_1_284);
	MAC_1_285: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_285, data_out=>output_MAC_1_285);
	MAC_1_286: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_286, data_out=>output_MAC_1_286);
	MAC_1_287: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_287, data_out=>output_MAC_1_287);
	MAC_1_288: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_288, data_out=>output_MAC_1_288);
	MAC_1_289: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_289, data_out=>output_MAC_1_289);
	MAC_1_290: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_290, data_out=>output_MAC_1_290);
	MAC_1_291: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_291, data_out=>output_MAC_1_291);
	MAC_1_292: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_292, data_out=>output_MAC_1_292);
	MAC_1_293: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_293, data_out=>output_MAC_1_293);
	MAC_1_294: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_294, data_out=>output_MAC_1_294);
	MAC_1_295: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_295, data_out=>output_MAC_1_295);
	MAC_1_296: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_296, data_out=>output_MAC_1_296);
	MAC_1_297: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_297, data_out=>output_MAC_1_297);
	MAC_1_298: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_298, data_out=>output_MAC_1_298);
	MAC_1_299: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_299, data_out=>output_MAC_1_299);
	MAC_1_300: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_300, data_out=>output_MAC_1_300);
	MAC_1_301: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_301, data_out=>output_MAC_1_301);
	MAC_1_302: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_302, data_out=>output_MAC_1_302);
	MAC_1_303: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_303, data_out=>output_MAC_1_303);
	MAC_1_304: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_304, data_out=>output_MAC_1_304);
	MAC_1_305: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_305, data_out=>output_MAC_1_305);
	MAC_1_306: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_306, data_out=>output_MAC_1_306);
	MAC_1_307: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_307, data_out=>output_MAC_1_307);
	MAC_1_308: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_308, data_out=>output_MAC_1_308);
	MAC_1_309: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_309, data_out=>output_MAC_1_309);
	MAC_1_310: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_310, data_out=>output_MAC_1_310);
	MAC_1_311: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_311, data_out=>output_MAC_1_311);
	MAC_1_312: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_312, data_out=>output_MAC_1_312);
	MAC_1_313: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_313, data_out=>output_MAC_1_313);
	MAC_1_314: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_314, data_out=>output_MAC_1_314);
	MAC_1_315: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_315, data_out=>output_MAC_1_315);
	MAC_1_316: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_316, data_out=>output_MAC_1_316);
	MAC_1_317: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_317, data_out=>output_MAC_1_317);
	MAC_1_318: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_318, data_out=>output_MAC_1_318);
	MAC_1_319: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_319, data_out=>output_MAC_1_319);
	MAC_1_320: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_320, data_out=>output_MAC_1_320);
	MAC_1_321: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_321, data_out=>output_MAC_1_321);
	MAC_1_322: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_322, data_out=>output_MAC_1_322);
	MAC_1_323: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_323, data_out=>output_MAC_1_323);
	MAC_1_324: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_324, data_out=>output_MAC_1_324);
	MAC_1_325: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_325, data_out=>output_MAC_1_325);
	MAC_1_326: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_326, data_out=>output_MAC_1_326);
	MAC_1_327: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_327, data_out=>output_MAC_1_327);
	MAC_1_328: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_328, data_out=>output_MAC_1_328);
	MAC_1_329: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_329, data_out=>output_MAC_1_329);
	MAC_1_330: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_330, data_out=>output_MAC_1_330);
	MAC_1_331: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_331, data_out=>output_MAC_1_331);
	MAC_1_332: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_332, data_out=>output_MAC_1_332);
	MAC_1_333: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_333, data_out=>output_MAC_1_333);
	MAC_1_334: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_334, data_out=>output_MAC_1_334);
	MAC_1_335: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_335, data_out=>output_MAC_1_335);
	MAC_1_336: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_336, data_out=>output_MAC_1_336);
	MAC_1_337: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_337, data_out=>output_MAC_1_337);
	MAC_1_338: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_338, data_out=>output_MAC_1_338);
	MAC_1_339: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_339, data_out=>output_MAC_1_339);
	MAC_1_340: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_340, data_out=>output_MAC_1_340);
	MAC_1_341: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_341, data_out=>output_MAC_1_341);
	MAC_1_342: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_342, data_out=>output_MAC_1_342);
	MAC_1_343: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_343, data_out=>output_MAC_1_343);
	MAC_1_344: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_344, data_out=>output_MAC_1_344);
	MAC_1_345: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_345, data_out=>output_MAC_1_345);
	MAC_1_346: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_346, data_out=>output_MAC_1_346);
	MAC_1_347: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_347, data_out=>output_MAC_1_347);
	MAC_1_348: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_348, data_out=>output_MAC_1_348);
	MAC_1_349: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_349, data_out=>output_MAC_1_349);
	MAC_1_350: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_350, data_out=>output_MAC_1_350);
	MAC_1_351: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_351, data_out=>output_MAC_1_351);
	MAC_1_352: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_352, data_out=>output_MAC_1_352);
	MAC_1_353: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_353, data_out=>output_MAC_1_353);
	MAC_1_354: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_354, data_out=>output_MAC_1_354);
	MAC_1_355: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_355, data_out=>output_MAC_1_355);
	MAC_1_356: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_356, data_out=>output_MAC_1_356);
	MAC_1_357: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_357, data_out=>output_MAC_1_357);
	MAC_1_358: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_358, data_out=>output_MAC_1_358);
	MAC_1_359: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_359, data_out=>output_MAC_1_359);
	MAC_1_360: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_360, data_out=>output_MAC_1_360);
	MAC_1_361: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_361, data_out=>output_MAC_1_361);
	MAC_1_362: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_362, data_out=>output_MAC_1_362);
	MAC_1_363: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_363, data_out=>output_MAC_1_363);
	MAC_1_364: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_364, data_out=>output_MAC_1_364);
	MAC_1_365: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_365, data_out=>output_MAC_1_365);
	MAC_1_366: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_366, data_out=>output_MAC_1_366);
	MAC_1_367: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_367, data_out=>output_MAC_1_367);
	MAC_1_368: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_368, data_out=>output_MAC_1_368);
	MAC_1_369: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_369, data_out=>output_MAC_1_369);
	MAC_1_370: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_370, data_out=>output_MAC_1_370);
	MAC_1_371: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_371, data_out=>output_MAC_1_371);
	MAC_1_372: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_372, data_out=>output_MAC_1_372);
	MAC_1_373: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_373, data_out=>output_MAC_1_373);
	MAC_1_374: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_374, data_out=>output_MAC_1_374);
	MAC_1_375: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_375, data_out=>output_MAC_1_375);
	MAC_1_376: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_376, data_out=>output_MAC_1_376);
	MAC_1_377: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_377, data_out=>output_MAC_1_377);
	MAC_1_378: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_378, data_out=>output_MAC_1_378);
	MAC_1_379: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_379, data_out=>output_MAC_1_379);
	MAC_1_380: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_380, data_out=>output_MAC_1_380);
	MAC_1_381: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_381, data_out=>output_MAC_1_381);
	MAC_1_382: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_382, data_out=>output_MAC_1_382);
	MAC_1_383: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_383, data_out=>output_MAC_1_383);
	MAC_1_384: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_384, data_out=>output_MAC_1_384);
	MAC_1_385: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_385, data_out=>output_MAC_1_385);
	MAC_1_386: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_386, data_out=>output_MAC_1_386);
	MAC_1_387: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_387, data_out=>output_MAC_1_387);
	MAC_1_388: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_388, data_out=>output_MAC_1_388);
	MAC_1_389: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_389, data_out=>output_MAC_1_389);
	MAC_1_390: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_390, data_out=>output_MAC_1_390);
	MAC_1_391: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_391, data_out=>output_MAC_1_391);
	MAC_1_392: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_392, data_out=>output_MAC_1_392);
	MAC_1_393: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_393, data_out=>output_MAC_1_393);
	MAC_1_394: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_394, data_out=>output_MAC_1_394);
	MAC_1_395: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_395, data_out=>output_MAC_1_395);
	MAC_1_396: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_396, data_out=>output_MAC_1_396);
	MAC_1_397: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_397, data_out=>output_MAC_1_397);
	MAC_1_398: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_398, data_out=>output_MAC_1_398);
	MAC_1_399: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_399, data_out=>output_MAC_1_399);
	MAC_1_400: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_400, data_out=>output_MAC_1_400);
	MAC_1_401: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_401, data_out=>output_MAC_1_401);
	MAC_1_402: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_402, data_out=>output_MAC_1_402);
	MAC_1_403: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_403, data_out=>output_MAC_1_403);
	MAC_1_404: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_404, data_out=>output_MAC_1_404);
	MAC_1_405: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_405, data_out=>output_MAC_1_405);
	MAC_1_406: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_406, data_out=>output_MAC_1_406);
	MAC_1_407: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_407, data_out=>output_MAC_1_407);
	MAC_1_408: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_408, data_out=>output_MAC_1_408);
	MAC_1_409: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_409, data_out=>output_MAC_1_409);
	MAC_1_410: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_410, data_out=>output_MAC_1_410);
	MAC_1_411: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_411, data_out=>output_MAC_1_411);
	MAC_1_412: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_412, data_out=>output_MAC_1_412);
	MAC_1_413: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_413, data_out=>output_MAC_1_413);
	MAC_1_414: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_414, data_out=>output_MAC_1_414);
	MAC_1_415: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_415, data_out=>output_MAC_1_415);
	MAC_1_416: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_416, data_out=>output_MAC_1_416);
	MAC_1_417: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_417, data_out=>output_MAC_1_417);
	MAC_1_418: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_418, data_out=>output_MAC_1_418);
	MAC_1_419: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_419, data_out=>output_MAC_1_419);
	MAC_1_420: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_420, data_out=>output_MAC_1_420);
	MAC_1_421: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_421, data_out=>output_MAC_1_421);
	MAC_1_422: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_422, data_out=>output_MAC_1_422);
	MAC_1_423: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_423, data_out=>output_MAC_1_423);
	MAC_1_424: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_424, data_out=>output_MAC_1_424);
	MAC_1_425: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_425, data_out=>output_MAC_1_425);
	MAC_1_426: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_426, data_out=>output_MAC_1_426);
	MAC_1_427: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_427, data_out=>output_MAC_1_427);
	MAC_1_428: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_428, data_out=>output_MAC_1_428);
	MAC_1_429: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_429, data_out=>output_MAC_1_429);
	MAC_1_430: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_430, data_out=>output_MAC_1_430);
	MAC_1_431: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_431, data_out=>output_MAC_1_431);
	MAC_1_432: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_432, data_out=>output_MAC_1_432);
	MAC_1_433: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_433, data_out=>output_MAC_1_433);
	MAC_1_434: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_434, data_out=>output_MAC_1_434);
	MAC_1_435: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_435, data_out=>output_MAC_1_435);
	MAC_1_436: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_436, data_out=>output_MAC_1_436);
	MAC_1_437: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_437, data_out=>output_MAC_1_437);
	MAC_1_438: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_438, data_out=>output_MAC_1_438);
	MAC_1_439: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_439, data_out=>output_MAC_1_439);
	MAC_1_440: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_440, data_out=>output_MAC_1_440);
	MAC_1_441: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_441, data_out=>output_MAC_1_441);
	MAC_1_442: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_442, data_out=>output_MAC_1_442);
	MAC_1_443: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_443, data_out=>output_MAC_1_443);
	MAC_1_444: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_444, data_out=>output_MAC_1_444);
	MAC_1_445: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_445, data_out=>output_MAC_1_445);
	MAC_1_446: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_446, data_out=>output_MAC_1_446);
	MAC_1_447: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_447, data_out=>output_MAC_1_447);
	MAC_1_448: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_448, data_out=>output_MAC_1_448);
	MAC_1_449: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_449, data_out=>output_MAC_1_449);
	MAC_1_450: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_450, data_out=>output_MAC_1_450);
	MAC_1_451: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_451, data_out=>output_MAC_1_451);
	MAC_1_452: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_452, data_out=>output_MAC_1_452);
	MAC_1_453: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_453, data_out=>output_MAC_1_453);
	MAC_1_454: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_454, data_out=>output_MAC_1_454);
	MAC_1_455: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_455, data_out=>output_MAC_1_455);
	MAC_1_456: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_456, data_out=>output_MAC_1_456);
	MAC_1_457: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_457, data_out=>output_MAC_1_457);
	MAC_1_458: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_458, data_out=>output_MAC_1_458);
	MAC_1_459: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_459, data_out=>output_MAC_1_459);
	MAC_1_460: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_460, data_out=>output_MAC_1_460);
	MAC_1_461: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_461, data_out=>output_MAC_1_461);
	MAC_1_462: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_462, data_out=>output_MAC_1_462);
	MAC_1_463: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_463, data_out=>output_MAC_1_463);
	MAC_1_464: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_464, data_out=>output_MAC_1_464);
	MAC_1_465: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_465, data_out=>output_MAC_1_465);
	MAC_1_466: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_466, data_out=>output_MAC_1_466);
	MAC_1_467: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_467, data_out=>output_MAC_1_467);
	MAC_1_468: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_468, data_out=>output_MAC_1_468);
	MAC_1_469: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_469, data_out=>output_MAC_1_469);
	MAC_1_470: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_470, data_out=>output_MAC_1_470);
	MAC_1_471: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_471, data_out=>output_MAC_1_471);
	MAC_1_472: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_472, data_out=>output_MAC_1_472);
	MAC_1_473: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_473, data_out=>output_MAC_1_473);
	MAC_1_474: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_474, data_out=>output_MAC_1_474);
	MAC_1_475: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_475, data_out=>output_MAC_1_475);
	MAC_1_476: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_476, data_out=>output_MAC_1_476);
	MAC_1_477: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_477, data_out=>output_MAC_1_477);
	MAC_1_478: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_478, data_out=>output_MAC_1_478);
	MAC_1_479: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_479, data_out=>output_MAC_1_479);
	MAC_1_480: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_480, data_out=>output_MAC_1_480);
	MAC_1_481: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_481, data_out=>output_MAC_1_481);
	MAC_1_482: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_482, data_out=>output_MAC_1_482);
	MAC_1_483: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_483, data_out=>output_MAC_1_483);
	MAC_1_484: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_484, data_out=>output_MAC_1_484);
	MAC_1_485: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_485, data_out=>output_MAC_1_485);
	MAC_1_486: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_486, data_out=>output_MAC_1_486);
	MAC_1_487: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_487, data_out=>output_MAC_1_487);
	MAC_1_488: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_488, data_out=>output_MAC_1_488);
	MAC_1_489: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_489, data_out=>output_MAC_1_489);
	MAC_1_490: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_490, data_out=>output_MAC_1_490);
	MAC_1_491: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_491, data_out=>output_MAC_1_491);
	MAC_1_492: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_492, data_out=>output_MAC_1_492);
	MAC_1_493: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_493, data_out=>output_MAC_1_493);
	MAC_1_494: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_494, data_out=>output_MAC_1_494);
	MAC_1_495: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_495, data_out=>output_MAC_1_495);
	MAC_1_496: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_496, data_out=>output_MAC_1_496);
	MAC_1_497: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_497, data_out=>output_MAC_1_497);
	MAC_1_498: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_498, data_out=>output_MAC_1_498);
	MAC_1_499: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_499, data_out=>output_MAC_1_499);
	MAC_1_500: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_500, data_out=>output_MAC_1_500);
	MAC_1_501: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_501, data_out=>output_MAC_1_501);
	MAC_1_502: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_502, data_out=>output_MAC_1_502);
	MAC_1_503: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_503, data_out=>output_MAC_1_503);
	MAC_1_504: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_504, data_out=>output_MAC_1_504);
	MAC_1_505: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_505, data_out=>output_MAC_1_505);
	MAC_1_506: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_506, data_out=>output_MAC_1_506);
	MAC_1_507: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_507, data_out=>output_MAC_1_507);
	MAC_1_508: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_508, data_out=>output_MAC_1_508);
	MAC_1_509: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_509, data_out=>output_MAC_1_509);
	MAC_1_510: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_510, data_out=>output_MAC_1_510);
	MAC_1_511: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_511, data_out=>output_MAC_1_511);
	MAC_1_512: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_512, data_out=>output_MAC_1_512);
	MAC_1_513: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_513, data_out=>output_MAC_1_513);
	MAC_1_514: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_514, data_out=>output_MAC_1_514);
	MAC_1_515: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_515, data_out=>output_MAC_1_515);
	MAC_1_516: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_516, data_out=>output_MAC_1_516);
	MAC_1_517: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_517, data_out=>output_MAC_1_517);
	MAC_1_518: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_518, data_out=>output_MAC_1_518);
	MAC_1_519: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_519, data_out=>output_MAC_1_519);
	MAC_1_520: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_520, data_out=>output_MAC_1_520);
	MAC_1_521: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_521, data_out=>output_MAC_1_521);
	MAC_1_522: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_522, data_out=>output_MAC_1_522);
	MAC_1_523: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_523, data_out=>output_MAC_1_523);
	MAC_1_524: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_524, data_out=>output_MAC_1_524);
	MAC_1_525: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_525, data_out=>output_MAC_1_525);
	MAC_1_526: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_526, data_out=>output_MAC_1_526);
	MAC_1_527: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_527, data_out=>output_MAC_1_527);
	MAC_1_528: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_528, data_out=>output_MAC_1_528);
	MAC_1_529: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_529, data_out=>output_MAC_1_529);
	MAC_1_530: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_530, data_out=>output_MAC_1_530);
	MAC_1_531: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_531, data_out=>output_MAC_1_531);
	MAC_1_532: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_532, data_out=>output_MAC_1_532);
	MAC_1_533: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_533, data_out=>output_MAC_1_533);
	MAC_1_534: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_534, data_out=>output_MAC_1_534);
	MAC_1_535: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_535, data_out=>output_MAC_1_535);
	MAC_1_536: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_536, data_out=>output_MAC_1_536);
	MAC_1_537: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_537, data_out=>output_MAC_1_537);
	MAC_1_538: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_538, data_out=>output_MAC_1_538);
	MAC_1_539: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_539, data_out=>output_MAC_1_539);
	MAC_1_540: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_540, data_out=>output_MAC_1_540);
	MAC_1_541: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_541, data_out=>output_MAC_1_541);
	MAC_1_542: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_542, data_out=>output_MAC_1_542);
	MAC_1_543: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_543, data_out=>output_MAC_1_543);
	MAC_1_544: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_544, data_out=>output_MAC_1_544);
	MAC_1_545: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_545, data_out=>output_MAC_1_545);
	MAC_1_546: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_546, data_out=>output_MAC_1_546);
	MAC_1_547: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_547, data_out=>output_MAC_1_547);
	MAC_1_548: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_548, data_out=>output_MAC_1_548);
	MAC_1_549: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_549, data_out=>output_MAC_1_549);
	MAC_1_550: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_550, data_out=>output_MAC_1_550);
	MAC_1_551: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_551, data_out=>output_MAC_1_551);
	MAC_1_552: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_552, data_out=>output_MAC_1_552);
	MAC_1_553: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_553, data_out=>output_MAC_1_553);
	MAC_1_554: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_554, data_out=>output_MAC_1_554);
	MAC_1_555: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_555, data_out=>output_MAC_1_555);
	MAC_1_556: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_556, data_out=>output_MAC_1_556);
	MAC_1_557: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_557, data_out=>output_MAC_1_557);
	MAC_1_558: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_558, data_out=>output_MAC_1_558);
	MAC_1_559: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_559, data_out=>output_MAC_1_559);
	MAC_1_560: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_560, data_out=>output_MAC_1_560);
	MAC_1_561: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_561, data_out=>output_MAC_1_561);
	MAC_1_562: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_562, data_out=>output_MAC_1_562);
	MAC_1_563: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_563, data_out=>output_MAC_1_563);
	MAC_1_564: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_564, data_out=>output_MAC_1_564);
	MAC_1_565: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_565, data_out=>output_MAC_1_565);
	MAC_1_566: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_566, data_out=>output_MAC_1_566);
	MAC_1_567: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_567, data_out=>output_MAC_1_567);
	MAC_1_568: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_568, data_out=>output_MAC_1_568);
	MAC_1_569: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_569, data_out=>output_MAC_1_569);
	MAC_1_570: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_570, data_out=>output_MAC_1_570);
	MAC_1_571: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_571, data_out=>output_MAC_1_571);
	MAC_1_572: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_572, data_out=>output_MAC_1_572);
	MAC_1_573: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_573, data_out=>output_MAC_1_573);
	MAC_1_574: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_574, data_out=>output_MAC_1_574);
	MAC_1_575: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_575, data_out=>output_MAC_1_575);
	MAC_1_576: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_576, data_out=>output_MAC_1_576);
	MAC_1_577: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_577, data_out=>output_MAC_1_577);
	MAC_1_578: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_578, data_out=>output_MAC_1_578);
	MAC_1_579: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_579, data_out=>output_MAC_1_579);
	MAC_1_580: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_580, data_out=>output_MAC_1_580);
	MAC_1_581: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_581, data_out=>output_MAC_1_581);
	MAC_1_582: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_582, data_out=>output_MAC_1_582);
	MAC_1_583: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_583, data_out=>output_MAC_1_583);
	MAC_1_584: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_584, data_out=>output_MAC_1_584);
	MAC_1_585: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_585, data_out=>output_MAC_1_585);
	MAC_1_586: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_586, data_out=>output_MAC_1_586);
	MAC_1_587: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_587, data_out=>output_MAC_1_587);
	MAC_1_588: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_588, data_out=>output_MAC_1_588);
	MAC_1_589: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_589, data_out=>output_MAC_1_589);
	MAC_1_590: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_590, data_out=>output_MAC_1_590);
	MAC_1_591: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_591, data_out=>output_MAC_1_591);
	MAC_1_592: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_592, data_out=>output_MAC_1_592);
	MAC_1_593: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_593, data_out=>output_MAC_1_593);
	MAC_1_594: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_594, data_out=>output_MAC_1_594);
	MAC_1_595: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_595, data_out=>output_MAC_1_595);
	MAC_1_596: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_596, data_out=>output_MAC_1_596);
	MAC_1_597: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_597, data_out=>output_MAC_1_597);
	MAC_1_598: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_598, data_out=>output_MAC_1_598);
	MAC_1_599: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_599, data_out=>output_MAC_1_599);
	MAC_1_600: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_600, data_out=>output_MAC_1_600);
	MAC_1_601: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_601, data_out=>output_MAC_1_601);
	MAC_1_602: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_602, data_out=>output_MAC_1_602);
	MAC_1_603: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_603, data_out=>output_MAC_1_603);
	MAC_1_604: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_604, data_out=>output_MAC_1_604);
	MAC_1_605: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_605, data_out=>output_MAC_1_605);
	MAC_1_606: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_606, data_out=>output_MAC_1_606);
	MAC_1_607: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_607, data_out=>output_MAC_1_607);
	MAC_1_608: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_608, data_out=>output_MAC_1_608);
	MAC_1_609: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_609, data_out=>output_MAC_1_609);
	MAC_1_610: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_610, data_out=>output_MAC_1_610);
	MAC_1_611: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_611, data_out=>output_MAC_1_611);
	MAC_1_612: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_612, data_out=>output_MAC_1_612);
	MAC_1_613: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_613, data_out=>output_MAC_1_613);
	MAC_1_614: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_614, data_out=>output_MAC_1_614);
	MAC_1_615: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_615, data_out=>output_MAC_1_615);
	MAC_1_616: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_616, data_out=>output_MAC_1_616);
	MAC_1_617: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_617, data_out=>output_MAC_1_617);
	MAC_1_618: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_618, data_out=>output_MAC_1_618);
	MAC_1_619: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_619, data_out=>output_MAC_1_619);
	MAC_1_620: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_620, data_out=>output_MAC_1_620);
	MAC_1_621: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_621, data_out=>output_MAC_1_621);
	MAC_1_622: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_622, data_out=>output_MAC_1_622);
	MAC_1_623: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_623, data_out=>output_MAC_1_623);
	MAC_1_624: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_624, data_out=>output_MAC_1_624);
	MAC_1_625: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_625, data_out=>output_MAC_1_625);
	MAC_1_626: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_626, data_out=>output_MAC_1_626);
	MAC_1_627: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_627, data_out=>output_MAC_1_627);
	MAC_1_628: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_628, data_out=>output_MAC_1_628);
	MAC_1_629: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_629, data_out=>output_MAC_1_629);
	MAC_1_630: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_630, data_out=>output_MAC_1_630);
	MAC_1_631: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_631, data_out=>output_MAC_1_631);
	MAC_1_632: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_632, data_out=>output_MAC_1_632);
	MAC_1_633: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_633, data_out=>output_MAC_1_633);
	MAC_1_634: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_634, data_out=>output_MAC_1_634);
	MAC_1_635: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_635, data_out=>output_MAC_1_635);
	MAC_1_636: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_636, data_out=>output_MAC_1_636);
	MAC_1_637: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_637, data_out=>output_MAC_1_637);
	MAC_1_638: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_638, data_out=>output_MAC_1_638);
	MAC_1_639: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_639, data_out=>output_MAC_1_639);
	MAC_1_640: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_640, data_out=>output_MAC_1_640);
	MAC_1_641: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_641, data_out=>output_MAC_1_641);
	MAC_1_642: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_642, data_out=>output_MAC_1_642);
	MAC_1_643: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_643, data_out=>output_MAC_1_643);
	MAC_1_644: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_644, data_out=>output_MAC_1_644);
	MAC_1_645: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_645, data_out=>output_MAC_1_645);
	MAC_1_646: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_646, data_out=>output_MAC_1_646);
	MAC_1_647: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_647, data_out=>output_MAC_1_647);
	MAC_1_648: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_648, data_out=>output_MAC_1_648);
	MAC_1_649: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_649, data_out=>output_MAC_1_649);
	MAC_1_650: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_650, data_out=>output_MAC_1_650);
	MAC_1_651: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_651, data_out=>output_MAC_1_651);
	MAC_1_652: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_652, data_out=>output_MAC_1_652);
	MAC_1_653: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_653, data_out=>output_MAC_1_653);
	MAC_1_654: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_654, data_out=>output_MAC_1_654);
	MAC_1_655: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_655, data_out=>output_MAC_1_655);
	MAC_1_656: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_656, data_out=>output_MAC_1_656);
	MAC_1_657: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_657, data_out=>output_MAC_1_657);
	MAC_1_658: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_658, data_out=>output_MAC_1_658);
	MAC_1_659: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_659, data_out=>output_MAC_1_659);
	MAC_1_660: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_660, data_out=>output_MAC_1_660);
	MAC_1_661: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_661, data_out=>output_MAC_1_661);
	MAC_1_662: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_662, data_out=>output_MAC_1_662);
	MAC_1_663: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_663, data_out=>output_MAC_1_663);
	MAC_1_664: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_664, data_out=>output_MAC_1_664);
	MAC_1_665: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_665, data_out=>output_MAC_1_665);
	MAC_1_666: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_666, data_out=>output_MAC_1_666);
	MAC_1_667: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_667, data_out=>output_MAC_1_667);
	MAC_1_668: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_668, data_out=>output_MAC_1_668);
	MAC_1_669: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_669, data_out=>output_MAC_1_669);
	MAC_1_670: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_670, data_out=>output_MAC_1_670);
	MAC_1_671: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_671, data_out=>output_MAC_1_671);
	MAC_1_672: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_672, data_out=>output_MAC_1_672);
	MAC_1_673: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_673, data_out=>output_MAC_1_673);
	MAC_1_674: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_674, data_out=>output_MAC_1_674);
	MAC_1_675: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_675, data_out=>output_MAC_1_675);
	MAC_1_676: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_676, data_out=>output_MAC_1_676);
	MAC_1_677: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_677, data_out=>output_MAC_1_677);
	MAC_1_678: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_678, data_out=>output_MAC_1_678);
	MAC_1_679: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_679, data_out=>output_MAC_1_679);
	MAC_1_680: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_680, data_out=>output_MAC_1_680);
	MAC_1_681: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_681, data_out=>output_MAC_1_681);
	MAC_1_682: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_682, data_out=>output_MAC_1_682);
	MAC_1_683: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_683, data_out=>output_MAC_1_683);
	MAC_1_684: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_684, data_out=>output_MAC_1_684);
	MAC_1_685: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_685, data_out=>output_MAC_1_685);
	MAC_1_686: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_686, data_out=>output_MAC_1_686);
	MAC_1_687: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_687, data_out=>output_MAC_1_687);
	MAC_1_688: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_688, data_out=>output_MAC_1_688);
	MAC_1_689: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_689, data_out=>output_MAC_1_689);
	MAC_1_690: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_690, data_out=>output_MAC_1_690);
	MAC_1_691: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_691, data_out=>output_MAC_1_691);
	MAC_1_692: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_692, data_out=>output_MAC_1_692);
	MAC_1_693: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_693, data_out=>output_MAC_1_693);
	MAC_1_694: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_694, data_out=>output_MAC_1_694);
	MAC_1_695: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_695, data_out=>output_MAC_1_695);
	MAC_1_696: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_696, data_out=>output_MAC_1_696);
	MAC_1_697: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_697, data_out=>output_MAC_1_697);
	MAC_1_698: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_698, data_out=>output_MAC_1_698);
	MAC_1_699: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_699, data_out=>output_MAC_1_699);
	MAC_1_700: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_700, data_out=>output_MAC_1_700);
	MAC_1_701: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_701, data_out=>output_MAC_1_701);
	MAC_1_702: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_702, data_out=>output_MAC_1_702);
	MAC_1_703: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_703, data_out=>output_MAC_1_703);
	MAC_1_704: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_704, data_out=>output_MAC_1_704);
	MAC_1_705: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_705, data_out=>output_MAC_1_705);
	MAC_1_706: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_706, data_out=>output_MAC_1_706);
	MAC_1_707: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_707, data_out=>output_MAC_1_707);
	MAC_1_708: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_708, data_out=>output_MAC_1_708);
	MAC_1_709: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_709, data_out=>output_MAC_1_709);
	MAC_1_710: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_710, data_out=>output_MAC_1_710);
	MAC_1_711: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_711, data_out=>output_MAC_1_711);
	MAC_1_712: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_712, data_out=>output_MAC_1_712);
	MAC_1_713: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_713, data_out=>output_MAC_1_713);
	MAC_1_714: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_714, data_out=>output_MAC_1_714);
	MAC_1_715: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_715, data_out=>output_MAC_1_715);
	MAC_1_716: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_716, data_out=>output_MAC_1_716);
	MAC_1_717: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_717, data_out=>output_MAC_1_717);
	MAC_1_718: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_718, data_out=>output_MAC_1_718);
	MAC_1_719: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_719, data_out=>output_MAC_1_719);
	MAC_1_720: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_720, data_out=>output_MAC_1_720);
	MAC_1_721: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_721, data_out=>output_MAC_1_721);
	MAC_1_722: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_722, data_out=>output_MAC_1_722);
	MAC_1_723: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_723, data_out=>output_MAC_1_723);
	MAC_1_724: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_724, data_out=>output_MAC_1_724);
	MAC_1_725: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_725, data_out=>output_MAC_1_725);
	MAC_1_726: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_726, data_out=>output_MAC_1_726);
	MAC_1_727: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_727, data_out=>output_MAC_1_727);
	MAC_1_728: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_728, data_out=>output_MAC_1_728);
	MAC_1_729: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_729, data_out=>output_MAC_1_729);
	MAC_1_730: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_730, data_out=>output_MAC_1_730);
	MAC_1_731: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_731, data_out=>output_MAC_1_731);
	MAC_1_732: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_732, data_out=>output_MAC_1_732);
	MAC_1_733: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_733, data_out=>output_MAC_1_733);
	MAC_1_734: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_734, data_out=>output_MAC_1_734);
	MAC_1_735: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_735, data_out=>output_MAC_1_735);
	MAC_1_736: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_736, data_out=>output_MAC_1_736);
	MAC_1_737: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_737, data_out=>output_MAC_1_737);
	MAC_1_738: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_738, data_out=>output_MAC_1_738);
	MAC_1_739: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_739, data_out=>output_MAC_1_739);
	MAC_1_740: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_740, data_out=>output_MAC_1_740);
	MAC_1_741: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_741, data_out=>output_MAC_1_741);
	MAC_1_742: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_742, data_out=>output_MAC_1_742);
	MAC_1_743: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_743, data_out=>output_MAC_1_743);
	MAC_1_744: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_744, data_out=>output_MAC_1_744);
	MAC_1_745: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_745, data_out=>output_MAC_1_745);
	MAC_1_746: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_746, data_out=>output_MAC_1_746);
	MAC_1_747: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_747, data_out=>output_MAC_1_747);
	MAC_1_748: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_748, data_out=>output_MAC_1_748);
	MAC_1_749: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_749, data_out=>output_MAC_1_749);
	MAC_1_750: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_750, data_out=>output_MAC_1_750);
	MAC_1_751: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_751, data_out=>output_MAC_1_751);
	MAC_1_752: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_752, data_out=>output_MAC_1_752);
	MAC_1_753: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_753, data_out=>output_MAC_1_753);
	MAC_1_754: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_754, data_out=>output_MAC_1_754);
	MAC_1_755: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_755, data_out=>output_MAC_1_755);
	MAC_1_756: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_756, data_out=>output_MAC_1_756);
	MAC_1_757: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_757, data_out=>output_MAC_1_757);
	MAC_1_758: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_758, data_out=>output_MAC_1_758);
	MAC_1_759: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_759, data_out=>output_MAC_1_759);
	MAC_1_760: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_760, data_out=>output_MAC_1_760);
	MAC_1_761: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_761, data_out=>output_MAC_1_761);
	MAC_1_762: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_762, data_out=>output_MAC_1_762);
	MAC_1_763: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_763, data_out=>output_MAC_1_763);
	MAC_1_764: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_764, data_out=>output_MAC_1_764);
	MAC_1_765: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_765, data_out=>output_MAC_1_765);
	MAC_1_766: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_766, data_out=>output_MAC_1_766);
	MAC_1_767: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_1, data_in_B=>input_col_767, data_out=>output_MAC_1_767);
	MAC_2_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_0, data_out=>output_MAC_2_0);
	MAC_2_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_1, data_out=>output_MAC_2_1);
	MAC_2_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_2, data_out=>output_MAC_2_2);
	MAC_2_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_3, data_out=>output_MAC_2_3);
	MAC_2_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_4, data_out=>output_MAC_2_4);
	MAC_2_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_5, data_out=>output_MAC_2_5);
	MAC_2_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_6, data_out=>output_MAC_2_6);
	MAC_2_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_7, data_out=>output_MAC_2_7);
	MAC_2_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_8, data_out=>output_MAC_2_8);
	MAC_2_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_9, data_out=>output_MAC_2_9);
	MAC_2_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_10, data_out=>output_MAC_2_10);
	MAC_2_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_11, data_out=>output_MAC_2_11);
	MAC_2_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_12, data_out=>output_MAC_2_12);
	MAC_2_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_13, data_out=>output_MAC_2_13);
	MAC_2_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_14, data_out=>output_MAC_2_14);
	MAC_2_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_15, data_out=>output_MAC_2_15);
	MAC_2_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_16, data_out=>output_MAC_2_16);
	MAC_2_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_17, data_out=>output_MAC_2_17);
	MAC_2_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_18, data_out=>output_MAC_2_18);
	MAC_2_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_19, data_out=>output_MAC_2_19);
	MAC_2_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_20, data_out=>output_MAC_2_20);
	MAC_2_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_21, data_out=>output_MAC_2_21);
	MAC_2_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_22, data_out=>output_MAC_2_22);
	MAC_2_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_23, data_out=>output_MAC_2_23);
	MAC_2_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_24, data_out=>output_MAC_2_24);
	MAC_2_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_25, data_out=>output_MAC_2_25);
	MAC_2_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_26, data_out=>output_MAC_2_26);
	MAC_2_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_27, data_out=>output_MAC_2_27);
	MAC_2_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_28, data_out=>output_MAC_2_28);
	MAC_2_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_29, data_out=>output_MAC_2_29);
	MAC_2_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_30, data_out=>output_MAC_2_30);
	MAC_2_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_31, data_out=>output_MAC_2_31);
	MAC_2_32: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_32, data_out=>output_MAC_2_32);
	MAC_2_33: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_33, data_out=>output_MAC_2_33);
	MAC_2_34: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_34, data_out=>output_MAC_2_34);
	MAC_2_35: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_35, data_out=>output_MAC_2_35);
	MAC_2_36: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_36, data_out=>output_MAC_2_36);
	MAC_2_37: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_37, data_out=>output_MAC_2_37);
	MAC_2_38: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_38, data_out=>output_MAC_2_38);
	MAC_2_39: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_39, data_out=>output_MAC_2_39);
	MAC_2_40: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_40, data_out=>output_MAC_2_40);
	MAC_2_41: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_41, data_out=>output_MAC_2_41);
	MAC_2_42: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_42, data_out=>output_MAC_2_42);
	MAC_2_43: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_43, data_out=>output_MAC_2_43);
	MAC_2_44: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_44, data_out=>output_MAC_2_44);
	MAC_2_45: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_45, data_out=>output_MAC_2_45);
	MAC_2_46: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_46, data_out=>output_MAC_2_46);
	MAC_2_47: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_47, data_out=>output_MAC_2_47);
	MAC_2_48: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_48, data_out=>output_MAC_2_48);
	MAC_2_49: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_49, data_out=>output_MAC_2_49);
	MAC_2_50: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_50, data_out=>output_MAC_2_50);
	MAC_2_51: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_51, data_out=>output_MAC_2_51);
	MAC_2_52: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_52, data_out=>output_MAC_2_52);
	MAC_2_53: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_53, data_out=>output_MAC_2_53);
	MAC_2_54: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_54, data_out=>output_MAC_2_54);
	MAC_2_55: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_55, data_out=>output_MAC_2_55);
	MAC_2_56: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_56, data_out=>output_MAC_2_56);
	MAC_2_57: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_57, data_out=>output_MAC_2_57);
	MAC_2_58: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_58, data_out=>output_MAC_2_58);
	MAC_2_59: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_59, data_out=>output_MAC_2_59);
	MAC_2_60: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_60, data_out=>output_MAC_2_60);
	MAC_2_61: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_61, data_out=>output_MAC_2_61);
	MAC_2_62: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_62, data_out=>output_MAC_2_62);
	MAC_2_63: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_63, data_out=>output_MAC_2_63);
	MAC_2_64: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_64, data_out=>output_MAC_2_64);
	MAC_2_65: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_65, data_out=>output_MAC_2_65);
	MAC_2_66: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_66, data_out=>output_MAC_2_66);
	MAC_2_67: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_67, data_out=>output_MAC_2_67);
	MAC_2_68: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_68, data_out=>output_MAC_2_68);
	MAC_2_69: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_69, data_out=>output_MAC_2_69);
	MAC_2_70: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_70, data_out=>output_MAC_2_70);
	MAC_2_71: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_71, data_out=>output_MAC_2_71);
	MAC_2_72: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_72, data_out=>output_MAC_2_72);
	MAC_2_73: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_73, data_out=>output_MAC_2_73);
	MAC_2_74: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_74, data_out=>output_MAC_2_74);
	MAC_2_75: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_75, data_out=>output_MAC_2_75);
	MAC_2_76: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_76, data_out=>output_MAC_2_76);
	MAC_2_77: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_77, data_out=>output_MAC_2_77);
	MAC_2_78: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_78, data_out=>output_MAC_2_78);
	MAC_2_79: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_79, data_out=>output_MAC_2_79);
	MAC_2_80: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_80, data_out=>output_MAC_2_80);
	MAC_2_81: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_81, data_out=>output_MAC_2_81);
	MAC_2_82: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_82, data_out=>output_MAC_2_82);
	MAC_2_83: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_83, data_out=>output_MAC_2_83);
	MAC_2_84: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_84, data_out=>output_MAC_2_84);
	MAC_2_85: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_85, data_out=>output_MAC_2_85);
	MAC_2_86: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_86, data_out=>output_MAC_2_86);
	MAC_2_87: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_87, data_out=>output_MAC_2_87);
	MAC_2_88: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_88, data_out=>output_MAC_2_88);
	MAC_2_89: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_89, data_out=>output_MAC_2_89);
	MAC_2_90: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_90, data_out=>output_MAC_2_90);
	MAC_2_91: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_91, data_out=>output_MAC_2_91);
	MAC_2_92: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_92, data_out=>output_MAC_2_92);
	MAC_2_93: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_93, data_out=>output_MAC_2_93);
	MAC_2_94: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_94, data_out=>output_MAC_2_94);
	MAC_2_95: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_95, data_out=>output_MAC_2_95);
	MAC_2_96: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_96, data_out=>output_MAC_2_96);
	MAC_2_97: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_97, data_out=>output_MAC_2_97);
	MAC_2_98: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_98, data_out=>output_MAC_2_98);
	MAC_2_99: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_99, data_out=>output_MAC_2_99);
	MAC_2_100: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_100, data_out=>output_MAC_2_100);
	MAC_2_101: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_101, data_out=>output_MAC_2_101);
	MAC_2_102: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_102, data_out=>output_MAC_2_102);
	MAC_2_103: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_103, data_out=>output_MAC_2_103);
	MAC_2_104: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_104, data_out=>output_MAC_2_104);
	MAC_2_105: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_105, data_out=>output_MAC_2_105);
	MAC_2_106: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_106, data_out=>output_MAC_2_106);
	MAC_2_107: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_107, data_out=>output_MAC_2_107);
	MAC_2_108: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_108, data_out=>output_MAC_2_108);
	MAC_2_109: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_109, data_out=>output_MAC_2_109);
	MAC_2_110: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_110, data_out=>output_MAC_2_110);
	MAC_2_111: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_111, data_out=>output_MAC_2_111);
	MAC_2_112: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_112, data_out=>output_MAC_2_112);
	MAC_2_113: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_113, data_out=>output_MAC_2_113);
	MAC_2_114: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_114, data_out=>output_MAC_2_114);
	MAC_2_115: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_115, data_out=>output_MAC_2_115);
	MAC_2_116: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_116, data_out=>output_MAC_2_116);
	MAC_2_117: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_117, data_out=>output_MAC_2_117);
	MAC_2_118: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_118, data_out=>output_MAC_2_118);
	MAC_2_119: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_119, data_out=>output_MAC_2_119);
	MAC_2_120: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_120, data_out=>output_MAC_2_120);
	MAC_2_121: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_121, data_out=>output_MAC_2_121);
	MAC_2_122: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_122, data_out=>output_MAC_2_122);
	MAC_2_123: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_123, data_out=>output_MAC_2_123);
	MAC_2_124: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_124, data_out=>output_MAC_2_124);
	MAC_2_125: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_125, data_out=>output_MAC_2_125);
	MAC_2_126: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_126, data_out=>output_MAC_2_126);
	MAC_2_127: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_127, data_out=>output_MAC_2_127);
	MAC_2_128: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_128, data_out=>output_MAC_2_128);
	MAC_2_129: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_129, data_out=>output_MAC_2_129);
	MAC_2_130: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_130, data_out=>output_MAC_2_130);
	MAC_2_131: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_131, data_out=>output_MAC_2_131);
	MAC_2_132: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_132, data_out=>output_MAC_2_132);
	MAC_2_133: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_133, data_out=>output_MAC_2_133);
	MAC_2_134: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_134, data_out=>output_MAC_2_134);
	MAC_2_135: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_135, data_out=>output_MAC_2_135);
	MAC_2_136: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_136, data_out=>output_MAC_2_136);
	MAC_2_137: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_137, data_out=>output_MAC_2_137);
	MAC_2_138: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_138, data_out=>output_MAC_2_138);
	MAC_2_139: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_139, data_out=>output_MAC_2_139);
	MAC_2_140: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_140, data_out=>output_MAC_2_140);
	MAC_2_141: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_141, data_out=>output_MAC_2_141);
	MAC_2_142: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_142, data_out=>output_MAC_2_142);
	MAC_2_143: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_143, data_out=>output_MAC_2_143);
	MAC_2_144: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_144, data_out=>output_MAC_2_144);
	MAC_2_145: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_145, data_out=>output_MAC_2_145);
	MAC_2_146: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_146, data_out=>output_MAC_2_146);
	MAC_2_147: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_147, data_out=>output_MAC_2_147);
	MAC_2_148: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_148, data_out=>output_MAC_2_148);
	MAC_2_149: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_149, data_out=>output_MAC_2_149);
	MAC_2_150: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_150, data_out=>output_MAC_2_150);
	MAC_2_151: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_151, data_out=>output_MAC_2_151);
	MAC_2_152: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_152, data_out=>output_MAC_2_152);
	MAC_2_153: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_153, data_out=>output_MAC_2_153);
	MAC_2_154: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_154, data_out=>output_MAC_2_154);
	MAC_2_155: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_155, data_out=>output_MAC_2_155);
	MAC_2_156: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_156, data_out=>output_MAC_2_156);
	MAC_2_157: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_157, data_out=>output_MAC_2_157);
	MAC_2_158: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_158, data_out=>output_MAC_2_158);
	MAC_2_159: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_159, data_out=>output_MAC_2_159);
	MAC_2_160: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_160, data_out=>output_MAC_2_160);
	MAC_2_161: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_161, data_out=>output_MAC_2_161);
	MAC_2_162: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_162, data_out=>output_MAC_2_162);
	MAC_2_163: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_163, data_out=>output_MAC_2_163);
	MAC_2_164: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_164, data_out=>output_MAC_2_164);
	MAC_2_165: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_165, data_out=>output_MAC_2_165);
	MAC_2_166: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_166, data_out=>output_MAC_2_166);
	MAC_2_167: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_167, data_out=>output_MAC_2_167);
	MAC_2_168: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_168, data_out=>output_MAC_2_168);
	MAC_2_169: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_169, data_out=>output_MAC_2_169);
	MAC_2_170: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_170, data_out=>output_MAC_2_170);
	MAC_2_171: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_171, data_out=>output_MAC_2_171);
	MAC_2_172: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_172, data_out=>output_MAC_2_172);
	MAC_2_173: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_173, data_out=>output_MAC_2_173);
	MAC_2_174: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_174, data_out=>output_MAC_2_174);
	MAC_2_175: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_175, data_out=>output_MAC_2_175);
	MAC_2_176: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_176, data_out=>output_MAC_2_176);
	MAC_2_177: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_177, data_out=>output_MAC_2_177);
	MAC_2_178: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_178, data_out=>output_MAC_2_178);
	MAC_2_179: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_179, data_out=>output_MAC_2_179);
	MAC_2_180: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_180, data_out=>output_MAC_2_180);
	MAC_2_181: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_181, data_out=>output_MAC_2_181);
	MAC_2_182: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_182, data_out=>output_MAC_2_182);
	MAC_2_183: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_183, data_out=>output_MAC_2_183);
	MAC_2_184: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_184, data_out=>output_MAC_2_184);
	MAC_2_185: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_185, data_out=>output_MAC_2_185);
	MAC_2_186: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_186, data_out=>output_MAC_2_186);
	MAC_2_187: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_187, data_out=>output_MAC_2_187);
	MAC_2_188: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_188, data_out=>output_MAC_2_188);
	MAC_2_189: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_189, data_out=>output_MAC_2_189);
	MAC_2_190: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_190, data_out=>output_MAC_2_190);
	MAC_2_191: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_191, data_out=>output_MAC_2_191);
	MAC_2_192: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_192, data_out=>output_MAC_2_192);
	MAC_2_193: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_193, data_out=>output_MAC_2_193);
	MAC_2_194: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_194, data_out=>output_MAC_2_194);
	MAC_2_195: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_195, data_out=>output_MAC_2_195);
	MAC_2_196: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_196, data_out=>output_MAC_2_196);
	MAC_2_197: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_197, data_out=>output_MAC_2_197);
	MAC_2_198: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_198, data_out=>output_MAC_2_198);
	MAC_2_199: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_199, data_out=>output_MAC_2_199);
	MAC_2_200: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_200, data_out=>output_MAC_2_200);
	MAC_2_201: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_201, data_out=>output_MAC_2_201);
	MAC_2_202: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_202, data_out=>output_MAC_2_202);
	MAC_2_203: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_203, data_out=>output_MAC_2_203);
	MAC_2_204: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_204, data_out=>output_MAC_2_204);
	MAC_2_205: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_205, data_out=>output_MAC_2_205);
	MAC_2_206: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_206, data_out=>output_MAC_2_206);
	MAC_2_207: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_207, data_out=>output_MAC_2_207);
	MAC_2_208: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_208, data_out=>output_MAC_2_208);
	MAC_2_209: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_209, data_out=>output_MAC_2_209);
	MAC_2_210: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_210, data_out=>output_MAC_2_210);
	MAC_2_211: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_211, data_out=>output_MAC_2_211);
	MAC_2_212: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_212, data_out=>output_MAC_2_212);
	MAC_2_213: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_213, data_out=>output_MAC_2_213);
	MAC_2_214: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_214, data_out=>output_MAC_2_214);
	MAC_2_215: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_215, data_out=>output_MAC_2_215);
	MAC_2_216: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_216, data_out=>output_MAC_2_216);
	MAC_2_217: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_217, data_out=>output_MAC_2_217);
	MAC_2_218: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_218, data_out=>output_MAC_2_218);
	MAC_2_219: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_219, data_out=>output_MAC_2_219);
	MAC_2_220: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_220, data_out=>output_MAC_2_220);
	MAC_2_221: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_221, data_out=>output_MAC_2_221);
	MAC_2_222: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_222, data_out=>output_MAC_2_222);
	MAC_2_223: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_223, data_out=>output_MAC_2_223);
	MAC_2_224: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_224, data_out=>output_MAC_2_224);
	MAC_2_225: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_225, data_out=>output_MAC_2_225);
	MAC_2_226: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_226, data_out=>output_MAC_2_226);
	MAC_2_227: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_227, data_out=>output_MAC_2_227);
	MAC_2_228: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_228, data_out=>output_MAC_2_228);
	MAC_2_229: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_229, data_out=>output_MAC_2_229);
	MAC_2_230: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_230, data_out=>output_MAC_2_230);
	MAC_2_231: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_231, data_out=>output_MAC_2_231);
	MAC_2_232: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_232, data_out=>output_MAC_2_232);
	MAC_2_233: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_233, data_out=>output_MAC_2_233);
	MAC_2_234: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_234, data_out=>output_MAC_2_234);
	MAC_2_235: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_235, data_out=>output_MAC_2_235);
	MAC_2_236: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_236, data_out=>output_MAC_2_236);
	MAC_2_237: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_237, data_out=>output_MAC_2_237);
	MAC_2_238: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_238, data_out=>output_MAC_2_238);
	MAC_2_239: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_239, data_out=>output_MAC_2_239);
	MAC_2_240: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_240, data_out=>output_MAC_2_240);
	MAC_2_241: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_241, data_out=>output_MAC_2_241);
	MAC_2_242: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_242, data_out=>output_MAC_2_242);
	MAC_2_243: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_243, data_out=>output_MAC_2_243);
	MAC_2_244: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_244, data_out=>output_MAC_2_244);
	MAC_2_245: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_245, data_out=>output_MAC_2_245);
	MAC_2_246: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_246, data_out=>output_MAC_2_246);
	MAC_2_247: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_247, data_out=>output_MAC_2_247);
	MAC_2_248: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_248, data_out=>output_MAC_2_248);
	MAC_2_249: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_249, data_out=>output_MAC_2_249);
	MAC_2_250: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_250, data_out=>output_MAC_2_250);
	MAC_2_251: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_251, data_out=>output_MAC_2_251);
	MAC_2_252: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_252, data_out=>output_MAC_2_252);
	MAC_2_253: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_253, data_out=>output_MAC_2_253);
	MAC_2_254: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_254, data_out=>output_MAC_2_254);
	MAC_2_255: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_255, data_out=>output_MAC_2_255);
	MAC_2_256: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_256, data_out=>output_MAC_2_256);
	MAC_2_257: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_257, data_out=>output_MAC_2_257);
	MAC_2_258: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_258, data_out=>output_MAC_2_258);
	MAC_2_259: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_259, data_out=>output_MAC_2_259);
	MAC_2_260: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_260, data_out=>output_MAC_2_260);
	MAC_2_261: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_261, data_out=>output_MAC_2_261);
	MAC_2_262: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_262, data_out=>output_MAC_2_262);
	MAC_2_263: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_263, data_out=>output_MAC_2_263);
	MAC_2_264: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_264, data_out=>output_MAC_2_264);
	MAC_2_265: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_265, data_out=>output_MAC_2_265);
	MAC_2_266: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_266, data_out=>output_MAC_2_266);
	MAC_2_267: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_267, data_out=>output_MAC_2_267);
	MAC_2_268: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_268, data_out=>output_MAC_2_268);
	MAC_2_269: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_269, data_out=>output_MAC_2_269);
	MAC_2_270: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_270, data_out=>output_MAC_2_270);
	MAC_2_271: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_271, data_out=>output_MAC_2_271);
	MAC_2_272: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_272, data_out=>output_MAC_2_272);
	MAC_2_273: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_273, data_out=>output_MAC_2_273);
	MAC_2_274: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_274, data_out=>output_MAC_2_274);
	MAC_2_275: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_275, data_out=>output_MAC_2_275);
	MAC_2_276: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_276, data_out=>output_MAC_2_276);
	MAC_2_277: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_277, data_out=>output_MAC_2_277);
	MAC_2_278: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_278, data_out=>output_MAC_2_278);
	MAC_2_279: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_279, data_out=>output_MAC_2_279);
	MAC_2_280: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_280, data_out=>output_MAC_2_280);
	MAC_2_281: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_281, data_out=>output_MAC_2_281);
	MAC_2_282: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_282, data_out=>output_MAC_2_282);
	MAC_2_283: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_283, data_out=>output_MAC_2_283);
	MAC_2_284: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_284, data_out=>output_MAC_2_284);
	MAC_2_285: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_285, data_out=>output_MAC_2_285);
	MAC_2_286: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_286, data_out=>output_MAC_2_286);
	MAC_2_287: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_287, data_out=>output_MAC_2_287);
	MAC_2_288: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_288, data_out=>output_MAC_2_288);
	MAC_2_289: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_289, data_out=>output_MAC_2_289);
	MAC_2_290: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_290, data_out=>output_MAC_2_290);
	MAC_2_291: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_291, data_out=>output_MAC_2_291);
	MAC_2_292: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_292, data_out=>output_MAC_2_292);
	MAC_2_293: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_293, data_out=>output_MAC_2_293);
	MAC_2_294: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_294, data_out=>output_MAC_2_294);
	MAC_2_295: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_295, data_out=>output_MAC_2_295);
	MAC_2_296: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_296, data_out=>output_MAC_2_296);
	MAC_2_297: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_297, data_out=>output_MAC_2_297);
	MAC_2_298: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_298, data_out=>output_MAC_2_298);
	MAC_2_299: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_299, data_out=>output_MAC_2_299);
	MAC_2_300: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_300, data_out=>output_MAC_2_300);
	MAC_2_301: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_301, data_out=>output_MAC_2_301);
	MAC_2_302: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_302, data_out=>output_MAC_2_302);
	MAC_2_303: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_303, data_out=>output_MAC_2_303);
	MAC_2_304: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_304, data_out=>output_MAC_2_304);
	MAC_2_305: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_305, data_out=>output_MAC_2_305);
	MAC_2_306: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_306, data_out=>output_MAC_2_306);
	MAC_2_307: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_307, data_out=>output_MAC_2_307);
	MAC_2_308: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_308, data_out=>output_MAC_2_308);
	MAC_2_309: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_309, data_out=>output_MAC_2_309);
	MAC_2_310: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_310, data_out=>output_MAC_2_310);
	MAC_2_311: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_311, data_out=>output_MAC_2_311);
	MAC_2_312: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_312, data_out=>output_MAC_2_312);
	MAC_2_313: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_313, data_out=>output_MAC_2_313);
	MAC_2_314: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_314, data_out=>output_MAC_2_314);
	MAC_2_315: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_315, data_out=>output_MAC_2_315);
	MAC_2_316: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_316, data_out=>output_MAC_2_316);
	MAC_2_317: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_317, data_out=>output_MAC_2_317);
	MAC_2_318: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_318, data_out=>output_MAC_2_318);
	MAC_2_319: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_319, data_out=>output_MAC_2_319);
	MAC_2_320: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_320, data_out=>output_MAC_2_320);
	MAC_2_321: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_321, data_out=>output_MAC_2_321);
	MAC_2_322: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_322, data_out=>output_MAC_2_322);
	MAC_2_323: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_323, data_out=>output_MAC_2_323);
	MAC_2_324: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_324, data_out=>output_MAC_2_324);
	MAC_2_325: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_325, data_out=>output_MAC_2_325);
	MAC_2_326: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_326, data_out=>output_MAC_2_326);
	MAC_2_327: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_327, data_out=>output_MAC_2_327);
	MAC_2_328: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_328, data_out=>output_MAC_2_328);
	MAC_2_329: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_329, data_out=>output_MAC_2_329);
	MAC_2_330: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_330, data_out=>output_MAC_2_330);
	MAC_2_331: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_331, data_out=>output_MAC_2_331);
	MAC_2_332: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_332, data_out=>output_MAC_2_332);
	MAC_2_333: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_333, data_out=>output_MAC_2_333);
	MAC_2_334: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_334, data_out=>output_MAC_2_334);
	MAC_2_335: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_335, data_out=>output_MAC_2_335);
	MAC_2_336: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_336, data_out=>output_MAC_2_336);
	MAC_2_337: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_337, data_out=>output_MAC_2_337);
	MAC_2_338: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_338, data_out=>output_MAC_2_338);
	MAC_2_339: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_339, data_out=>output_MAC_2_339);
	MAC_2_340: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_340, data_out=>output_MAC_2_340);
	MAC_2_341: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_341, data_out=>output_MAC_2_341);
	MAC_2_342: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_342, data_out=>output_MAC_2_342);
	MAC_2_343: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_343, data_out=>output_MAC_2_343);
	MAC_2_344: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_344, data_out=>output_MAC_2_344);
	MAC_2_345: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_345, data_out=>output_MAC_2_345);
	MAC_2_346: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_346, data_out=>output_MAC_2_346);
	MAC_2_347: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_347, data_out=>output_MAC_2_347);
	MAC_2_348: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_348, data_out=>output_MAC_2_348);
	MAC_2_349: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_349, data_out=>output_MAC_2_349);
	MAC_2_350: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_350, data_out=>output_MAC_2_350);
	MAC_2_351: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_351, data_out=>output_MAC_2_351);
	MAC_2_352: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_352, data_out=>output_MAC_2_352);
	MAC_2_353: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_353, data_out=>output_MAC_2_353);
	MAC_2_354: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_354, data_out=>output_MAC_2_354);
	MAC_2_355: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_355, data_out=>output_MAC_2_355);
	MAC_2_356: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_356, data_out=>output_MAC_2_356);
	MAC_2_357: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_357, data_out=>output_MAC_2_357);
	MAC_2_358: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_358, data_out=>output_MAC_2_358);
	MAC_2_359: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_359, data_out=>output_MAC_2_359);
	MAC_2_360: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_360, data_out=>output_MAC_2_360);
	MAC_2_361: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_361, data_out=>output_MAC_2_361);
	MAC_2_362: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_362, data_out=>output_MAC_2_362);
	MAC_2_363: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_363, data_out=>output_MAC_2_363);
	MAC_2_364: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_364, data_out=>output_MAC_2_364);
	MAC_2_365: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_365, data_out=>output_MAC_2_365);
	MAC_2_366: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_366, data_out=>output_MAC_2_366);
	MAC_2_367: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_367, data_out=>output_MAC_2_367);
	MAC_2_368: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_368, data_out=>output_MAC_2_368);
	MAC_2_369: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_369, data_out=>output_MAC_2_369);
	MAC_2_370: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_370, data_out=>output_MAC_2_370);
	MAC_2_371: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_371, data_out=>output_MAC_2_371);
	MAC_2_372: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_372, data_out=>output_MAC_2_372);
	MAC_2_373: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_373, data_out=>output_MAC_2_373);
	MAC_2_374: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_374, data_out=>output_MAC_2_374);
	MAC_2_375: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_375, data_out=>output_MAC_2_375);
	MAC_2_376: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_376, data_out=>output_MAC_2_376);
	MAC_2_377: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_377, data_out=>output_MAC_2_377);
	MAC_2_378: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_378, data_out=>output_MAC_2_378);
	MAC_2_379: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_379, data_out=>output_MAC_2_379);
	MAC_2_380: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_380, data_out=>output_MAC_2_380);
	MAC_2_381: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_381, data_out=>output_MAC_2_381);
	MAC_2_382: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_382, data_out=>output_MAC_2_382);
	MAC_2_383: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_383, data_out=>output_MAC_2_383);
	MAC_2_384: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_384, data_out=>output_MAC_2_384);
	MAC_2_385: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_385, data_out=>output_MAC_2_385);
	MAC_2_386: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_386, data_out=>output_MAC_2_386);
	MAC_2_387: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_387, data_out=>output_MAC_2_387);
	MAC_2_388: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_388, data_out=>output_MAC_2_388);
	MAC_2_389: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_389, data_out=>output_MAC_2_389);
	MAC_2_390: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_390, data_out=>output_MAC_2_390);
	MAC_2_391: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_391, data_out=>output_MAC_2_391);
	MAC_2_392: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_392, data_out=>output_MAC_2_392);
	MAC_2_393: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_393, data_out=>output_MAC_2_393);
	MAC_2_394: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_394, data_out=>output_MAC_2_394);
	MAC_2_395: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_395, data_out=>output_MAC_2_395);
	MAC_2_396: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_396, data_out=>output_MAC_2_396);
	MAC_2_397: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_397, data_out=>output_MAC_2_397);
	MAC_2_398: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_398, data_out=>output_MAC_2_398);
	MAC_2_399: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_399, data_out=>output_MAC_2_399);
	MAC_2_400: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_400, data_out=>output_MAC_2_400);
	MAC_2_401: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_401, data_out=>output_MAC_2_401);
	MAC_2_402: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_402, data_out=>output_MAC_2_402);
	MAC_2_403: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_403, data_out=>output_MAC_2_403);
	MAC_2_404: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_404, data_out=>output_MAC_2_404);
	MAC_2_405: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_405, data_out=>output_MAC_2_405);
	MAC_2_406: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_406, data_out=>output_MAC_2_406);
	MAC_2_407: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_407, data_out=>output_MAC_2_407);
	MAC_2_408: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_408, data_out=>output_MAC_2_408);
	MAC_2_409: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_409, data_out=>output_MAC_2_409);
	MAC_2_410: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_410, data_out=>output_MAC_2_410);
	MAC_2_411: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_411, data_out=>output_MAC_2_411);
	MAC_2_412: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_412, data_out=>output_MAC_2_412);
	MAC_2_413: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_413, data_out=>output_MAC_2_413);
	MAC_2_414: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_414, data_out=>output_MAC_2_414);
	MAC_2_415: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_415, data_out=>output_MAC_2_415);
	MAC_2_416: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_416, data_out=>output_MAC_2_416);
	MAC_2_417: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_417, data_out=>output_MAC_2_417);
	MAC_2_418: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_418, data_out=>output_MAC_2_418);
	MAC_2_419: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_419, data_out=>output_MAC_2_419);
	MAC_2_420: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_420, data_out=>output_MAC_2_420);
	MAC_2_421: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_421, data_out=>output_MAC_2_421);
	MAC_2_422: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_422, data_out=>output_MAC_2_422);
	MAC_2_423: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_423, data_out=>output_MAC_2_423);
	MAC_2_424: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_424, data_out=>output_MAC_2_424);
	MAC_2_425: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_425, data_out=>output_MAC_2_425);
	MAC_2_426: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_426, data_out=>output_MAC_2_426);
	MAC_2_427: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_427, data_out=>output_MAC_2_427);
	MAC_2_428: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_428, data_out=>output_MAC_2_428);
	MAC_2_429: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_429, data_out=>output_MAC_2_429);
	MAC_2_430: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_430, data_out=>output_MAC_2_430);
	MAC_2_431: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_431, data_out=>output_MAC_2_431);
	MAC_2_432: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_432, data_out=>output_MAC_2_432);
	MAC_2_433: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_433, data_out=>output_MAC_2_433);
	MAC_2_434: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_434, data_out=>output_MAC_2_434);
	MAC_2_435: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_435, data_out=>output_MAC_2_435);
	MAC_2_436: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_436, data_out=>output_MAC_2_436);
	MAC_2_437: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_437, data_out=>output_MAC_2_437);
	MAC_2_438: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_438, data_out=>output_MAC_2_438);
	MAC_2_439: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_439, data_out=>output_MAC_2_439);
	MAC_2_440: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_440, data_out=>output_MAC_2_440);
	MAC_2_441: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_441, data_out=>output_MAC_2_441);
	MAC_2_442: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_442, data_out=>output_MAC_2_442);
	MAC_2_443: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_443, data_out=>output_MAC_2_443);
	MAC_2_444: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_444, data_out=>output_MAC_2_444);
	MAC_2_445: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_445, data_out=>output_MAC_2_445);
	MAC_2_446: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_446, data_out=>output_MAC_2_446);
	MAC_2_447: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_447, data_out=>output_MAC_2_447);
	MAC_2_448: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_448, data_out=>output_MAC_2_448);
	MAC_2_449: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_449, data_out=>output_MAC_2_449);
	MAC_2_450: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_450, data_out=>output_MAC_2_450);
	MAC_2_451: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_451, data_out=>output_MAC_2_451);
	MAC_2_452: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_452, data_out=>output_MAC_2_452);
	MAC_2_453: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_453, data_out=>output_MAC_2_453);
	MAC_2_454: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_454, data_out=>output_MAC_2_454);
	MAC_2_455: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_455, data_out=>output_MAC_2_455);
	MAC_2_456: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_456, data_out=>output_MAC_2_456);
	MAC_2_457: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_457, data_out=>output_MAC_2_457);
	MAC_2_458: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_458, data_out=>output_MAC_2_458);
	MAC_2_459: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_459, data_out=>output_MAC_2_459);
	MAC_2_460: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_460, data_out=>output_MAC_2_460);
	MAC_2_461: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_461, data_out=>output_MAC_2_461);
	MAC_2_462: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_462, data_out=>output_MAC_2_462);
	MAC_2_463: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_463, data_out=>output_MAC_2_463);
	MAC_2_464: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_464, data_out=>output_MAC_2_464);
	MAC_2_465: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_465, data_out=>output_MAC_2_465);
	MAC_2_466: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_466, data_out=>output_MAC_2_466);
	MAC_2_467: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_467, data_out=>output_MAC_2_467);
	MAC_2_468: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_468, data_out=>output_MAC_2_468);
	MAC_2_469: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_469, data_out=>output_MAC_2_469);
	MAC_2_470: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_470, data_out=>output_MAC_2_470);
	MAC_2_471: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_471, data_out=>output_MAC_2_471);
	MAC_2_472: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_472, data_out=>output_MAC_2_472);
	MAC_2_473: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_473, data_out=>output_MAC_2_473);
	MAC_2_474: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_474, data_out=>output_MAC_2_474);
	MAC_2_475: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_475, data_out=>output_MAC_2_475);
	MAC_2_476: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_476, data_out=>output_MAC_2_476);
	MAC_2_477: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_477, data_out=>output_MAC_2_477);
	MAC_2_478: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_478, data_out=>output_MAC_2_478);
	MAC_2_479: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_479, data_out=>output_MAC_2_479);
	MAC_2_480: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_480, data_out=>output_MAC_2_480);
	MAC_2_481: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_481, data_out=>output_MAC_2_481);
	MAC_2_482: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_482, data_out=>output_MAC_2_482);
	MAC_2_483: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_483, data_out=>output_MAC_2_483);
	MAC_2_484: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_484, data_out=>output_MAC_2_484);
	MAC_2_485: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_485, data_out=>output_MAC_2_485);
	MAC_2_486: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_486, data_out=>output_MAC_2_486);
	MAC_2_487: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_487, data_out=>output_MAC_2_487);
	MAC_2_488: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_488, data_out=>output_MAC_2_488);
	MAC_2_489: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_489, data_out=>output_MAC_2_489);
	MAC_2_490: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_490, data_out=>output_MAC_2_490);
	MAC_2_491: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_491, data_out=>output_MAC_2_491);
	MAC_2_492: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_492, data_out=>output_MAC_2_492);
	MAC_2_493: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_493, data_out=>output_MAC_2_493);
	MAC_2_494: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_494, data_out=>output_MAC_2_494);
	MAC_2_495: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_495, data_out=>output_MAC_2_495);
	MAC_2_496: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_496, data_out=>output_MAC_2_496);
	MAC_2_497: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_497, data_out=>output_MAC_2_497);
	MAC_2_498: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_498, data_out=>output_MAC_2_498);
	MAC_2_499: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_499, data_out=>output_MAC_2_499);
	MAC_2_500: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_500, data_out=>output_MAC_2_500);
	MAC_2_501: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_501, data_out=>output_MAC_2_501);
	MAC_2_502: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_502, data_out=>output_MAC_2_502);
	MAC_2_503: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_503, data_out=>output_MAC_2_503);
	MAC_2_504: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_504, data_out=>output_MAC_2_504);
	MAC_2_505: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_505, data_out=>output_MAC_2_505);
	MAC_2_506: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_506, data_out=>output_MAC_2_506);
	MAC_2_507: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_507, data_out=>output_MAC_2_507);
	MAC_2_508: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_508, data_out=>output_MAC_2_508);
	MAC_2_509: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_509, data_out=>output_MAC_2_509);
	MAC_2_510: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_510, data_out=>output_MAC_2_510);
	MAC_2_511: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_511, data_out=>output_MAC_2_511);
	MAC_2_512: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_512, data_out=>output_MAC_2_512);
	MAC_2_513: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_513, data_out=>output_MAC_2_513);
	MAC_2_514: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_514, data_out=>output_MAC_2_514);
	MAC_2_515: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_515, data_out=>output_MAC_2_515);
	MAC_2_516: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_516, data_out=>output_MAC_2_516);
	MAC_2_517: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_517, data_out=>output_MAC_2_517);
	MAC_2_518: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_518, data_out=>output_MAC_2_518);
	MAC_2_519: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_519, data_out=>output_MAC_2_519);
	MAC_2_520: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_520, data_out=>output_MAC_2_520);
	MAC_2_521: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_521, data_out=>output_MAC_2_521);
	MAC_2_522: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_522, data_out=>output_MAC_2_522);
	MAC_2_523: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_523, data_out=>output_MAC_2_523);
	MAC_2_524: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_524, data_out=>output_MAC_2_524);
	MAC_2_525: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_525, data_out=>output_MAC_2_525);
	MAC_2_526: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_526, data_out=>output_MAC_2_526);
	MAC_2_527: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_527, data_out=>output_MAC_2_527);
	MAC_2_528: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_528, data_out=>output_MAC_2_528);
	MAC_2_529: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_529, data_out=>output_MAC_2_529);
	MAC_2_530: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_530, data_out=>output_MAC_2_530);
	MAC_2_531: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_531, data_out=>output_MAC_2_531);
	MAC_2_532: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_532, data_out=>output_MAC_2_532);
	MAC_2_533: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_533, data_out=>output_MAC_2_533);
	MAC_2_534: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_534, data_out=>output_MAC_2_534);
	MAC_2_535: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_535, data_out=>output_MAC_2_535);
	MAC_2_536: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_536, data_out=>output_MAC_2_536);
	MAC_2_537: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_537, data_out=>output_MAC_2_537);
	MAC_2_538: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_538, data_out=>output_MAC_2_538);
	MAC_2_539: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_539, data_out=>output_MAC_2_539);
	MAC_2_540: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_540, data_out=>output_MAC_2_540);
	MAC_2_541: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_541, data_out=>output_MAC_2_541);
	MAC_2_542: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_542, data_out=>output_MAC_2_542);
	MAC_2_543: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_543, data_out=>output_MAC_2_543);
	MAC_2_544: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_544, data_out=>output_MAC_2_544);
	MAC_2_545: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_545, data_out=>output_MAC_2_545);
	MAC_2_546: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_546, data_out=>output_MAC_2_546);
	MAC_2_547: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_547, data_out=>output_MAC_2_547);
	MAC_2_548: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_548, data_out=>output_MAC_2_548);
	MAC_2_549: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_549, data_out=>output_MAC_2_549);
	MAC_2_550: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_550, data_out=>output_MAC_2_550);
	MAC_2_551: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_551, data_out=>output_MAC_2_551);
	MAC_2_552: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_552, data_out=>output_MAC_2_552);
	MAC_2_553: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_553, data_out=>output_MAC_2_553);
	MAC_2_554: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_554, data_out=>output_MAC_2_554);
	MAC_2_555: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_555, data_out=>output_MAC_2_555);
	MAC_2_556: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_556, data_out=>output_MAC_2_556);
	MAC_2_557: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_557, data_out=>output_MAC_2_557);
	MAC_2_558: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_558, data_out=>output_MAC_2_558);
	MAC_2_559: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_559, data_out=>output_MAC_2_559);
	MAC_2_560: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_560, data_out=>output_MAC_2_560);
	MAC_2_561: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_561, data_out=>output_MAC_2_561);
	MAC_2_562: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_562, data_out=>output_MAC_2_562);
	MAC_2_563: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_563, data_out=>output_MAC_2_563);
	MAC_2_564: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_564, data_out=>output_MAC_2_564);
	MAC_2_565: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_565, data_out=>output_MAC_2_565);
	MAC_2_566: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_566, data_out=>output_MAC_2_566);
	MAC_2_567: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_567, data_out=>output_MAC_2_567);
	MAC_2_568: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_568, data_out=>output_MAC_2_568);
	MAC_2_569: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_569, data_out=>output_MAC_2_569);
	MAC_2_570: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_570, data_out=>output_MAC_2_570);
	MAC_2_571: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_571, data_out=>output_MAC_2_571);
	MAC_2_572: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_572, data_out=>output_MAC_2_572);
	MAC_2_573: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_573, data_out=>output_MAC_2_573);
	MAC_2_574: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_574, data_out=>output_MAC_2_574);
	MAC_2_575: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_575, data_out=>output_MAC_2_575);
	MAC_2_576: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_576, data_out=>output_MAC_2_576);
	MAC_2_577: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_577, data_out=>output_MAC_2_577);
	MAC_2_578: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_578, data_out=>output_MAC_2_578);
	MAC_2_579: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_579, data_out=>output_MAC_2_579);
	MAC_2_580: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_580, data_out=>output_MAC_2_580);
	MAC_2_581: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_581, data_out=>output_MAC_2_581);
	MAC_2_582: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_582, data_out=>output_MAC_2_582);
	MAC_2_583: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_583, data_out=>output_MAC_2_583);
	MAC_2_584: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_584, data_out=>output_MAC_2_584);
	MAC_2_585: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_585, data_out=>output_MAC_2_585);
	MAC_2_586: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_586, data_out=>output_MAC_2_586);
	MAC_2_587: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_587, data_out=>output_MAC_2_587);
	MAC_2_588: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_588, data_out=>output_MAC_2_588);
	MAC_2_589: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_589, data_out=>output_MAC_2_589);
	MAC_2_590: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_590, data_out=>output_MAC_2_590);
	MAC_2_591: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_591, data_out=>output_MAC_2_591);
	MAC_2_592: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_592, data_out=>output_MAC_2_592);
	MAC_2_593: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_593, data_out=>output_MAC_2_593);
	MAC_2_594: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_594, data_out=>output_MAC_2_594);
	MAC_2_595: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_595, data_out=>output_MAC_2_595);
	MAC_2_596: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_596, data_out=>output_MAC_2_596);
	MAC_2_597: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_597, data_out=>output_MAC_2_597);
	MAC_2_598: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_598, data_out=>output_MAC_2_598);
	MAC_2_599: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_599, data_out=>output_MAC_2_599);
	MAC_2_600: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_600, data_out=>output_MAC_2_600);
	MAC_2_601: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_601, data_out=>output_MAC_2_601);
	MAC_2_602: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_602, data_out=>output_MAC_2_602);
	MAC_2_603: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_603, data_out=>output_MAC_2_603);
	MAC_2_604: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_604, data_out=>output_MAC_2_604);
	MAC_2_605: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_605, data_out=>output_MAC_2_605);
	MAC_2_606: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_606, data_out=>output_MAC_2_606);
	MAC_2_607: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_607, data_out=>output_MAC_2_607);
	MAC_2_608: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_608, data_out=>output_MAC_2_608);
	MAC_2_609: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_609, data_out=>output_MAC_2_609);
	MAC_2_610: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_610, data_out=>output_MAC_2_610);
	MAC_2_611: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_611, data_out=>output_MAC_2_611);
	MAC_2_612: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_612, data_out=>output_MAC_2_612);
	MAC_2_613: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_613, data_out=>output_MAC_2_613);
	MAC_2_614: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_614, data_out=>output_MAC_2_614);
	MAC_2_615: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_615, data_out=>output_MAC_2_615);
	MAC_2_616: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_616, data_out=>output_MAC_2_616);
	MAC_2_617: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_617, data_out=>output_MAC_2_617);
	MAC_2_618: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_618, data_out=>output_MAC_2_618);
	MAC_2_619: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_619, data_out=>output_MAC_2_619);
	MAC_2_620: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_620, data_out=>output_MAC_2_620);
	MAC_2_621: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_621, data_out=>output_MAC_2_621);
	MAC_2_622: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_622, data_out=>output_MAC_2_622);
	MAC_2_623: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_623, data_out=>output_MAC_2_623);
	MAC_2_624: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_624, data_out=>output_MAC_2_624);
	MAC_2_625: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_625, data_out=>output_MAC_2_625);
	MAC_2_626: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_626, data_out=>output_MAC_2_626);
	MAC_2_627: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_627, data_out=>output_MAC_2_627);
	MAC_2_628: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_628, data_out=>output_MAC_2_628);
	MAC_2_629: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_629, data_out=>output_MAC_2_629);
	MAC_2_630: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_630, data_out=>output_MAC_2_630);
	MAC_2_631: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_631, data_out=>output_MAC_2_631);
	MAC_2_632: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_632, data_out=>output_MAC_2_632);
	MAC_2_633: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_633, data_out=>output_MAC_2_633);
	MAC_2_634: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_634, data_out=>output_MAC_2_634);
	MAC_2_635: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_635, data_out=>output_MAC_2_635);
	MAC_2_636: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_636, data_out=>output_MAC_2_636);
	MAC_2_637: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_637, data_out=>output_MAC_2_637);
	MAC_2_638: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_638, data_out=>output_MAC_2_638);
	MAC_2_639: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_639, data_out=>output_MAC_2_639);
	MAC_2_640: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_640, data_out=>output_MAC_2_640);
	MAC_2_641: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_641, data_out=>output_MAC_2_641);
	MAC_2_642: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_642, data_out=>output_MAC_2_642);
	MAC_2_643: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_643, data_out=>output_MAC_2_643);
	MAC_2_644: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_644, data_out=>output_MAC_2_644);
	MAC_2_645: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_645, data_out=>output_MAC_2_645);
	MAC_2_646: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_646, data_out=>output_MAC_2_646);
	MAC_2_647: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_647, data_out=>output_MAC_2_647);
	MAC_2_648: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_648, data_out=>output_MAC_2_648);
	MAC_2_649: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_649, data_out=>output_MAC_2_649);
	MAC_2_650: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_650, data_out=>output_MAC_2_650);
	MAC_2_651: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_651, data_out=>output_MAC_2_651);
	MAC_2_652: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_652, data_out=>output_MAC_2_652);
	MAC_2_653: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_653, data_out=>output_MAC_2_653);
	MAC_2_654: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_654, data_out=>output_MAC_2_654);
	MAC_2_655: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_655, data_out=>output_MAC_2_655);
	MAC_2_656: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_656, data_out=>output_MAC_2_656);
	MAC_2_657: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_657, data_out=>output_MAC_2_657);
	MAC_2_658: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_658, data_out=>output_MAC_2_658);
	MAC_2_659: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_659, data_out=>output_MAC_2_659);
	MAC_2_660: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_660, data_out=>output_MAC_2_660);
	MAC_2_661: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_661, data_out=>output_MAC_2_661);
	MAC_2_662: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_662, data_out=>output_MAC_2_662);
	MAC_2_663: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_663, data_out=>output_MAC_2_663);
	MAC_2_664: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_664, data_out=>output_MAC_2_664);
	MAC_2_665: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_665, data_out=>output_MAC_2_665);
	MAC_2_666: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_666, data_out=>output_MAC_2_666);
	MAC_2_667: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_667, data_out=>output_MAC_2_667);
	MAC_2_668: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_668, data_out=>output_MAC_2_668);
	MAC_2_669: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_669, data_out=>output_MAC_2_669);
	MAC_2_670: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_670, data_out=>output_MAC_2_670);
	MAC_2_671: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_671, data_out=>output_MAC_2_671);
	MAC_2_672: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_672, data_out=>output_MAC_2_672);
	MAC_2_673: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_673, data_out=>output_MAC_2_673);
	MAC_2_674: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_674, data_out=>output_MAC_2_674);
	MAC_2_675: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_675, data_out=>output_MAC_2_675);
	MAC_2_676: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_676, data_out=>output_MAC_2_676);
	MAC_2_677: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_677, data_out=>output_MAC_2_677);
	MAC_2_678: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_678, data_out=>output_MAC_2_678);
	MAC_2_679: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_679, data_out=>output_MAC_2_679);
	MAC_2_680: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_680, data_out=>output_MAC_2_680);
	MAC_2_681: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_681, data_out=>output_MAC_2_681);
	MAC_2_682: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_682, data_out=>output_MAC_2_682);
	MAC_2_683: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_683, data_out=>output_MAC_2_683);
	MAC_2_684: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_684, data_out=>output_MAC_2_684);
	MAC_2_685: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_685, data_out=>output_MAC_2_685);
	MAC_2_686: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_686, data_out=>output_MAC_2_686);
	MAC_2_687: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_687, data_out=>output_MAC_2_687);
	MAC_2_688: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_688, data_out=>output_MAC_2_688);
	MAC_2_689: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_689, data_out=>output_MAC_2_689);
	MAC_2_690: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_690, data_out=>output_MAC_2_690);
	MAC_2_691: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_691, data_out=>output_MAC_2_691);
	MAC_2_692: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_692, data_out=>output_MAC_2_692);
	MAC_2_693: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_693, data_out=>output_MAC_2_693);
	MAC_2_694: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_694, data_out=>output_MAC_2_694);
	MAC_2_695: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_695, data_out=>output_MAC_2_695);
	MAC_2_696: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_696, data_out=>output_MAC_2_696);
	MAC_2_697: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_697, data_out=>output_MAC_2_697);
	MAC_2_698: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_698, data_out=>output_MAC_2_698);
	MAC_2_699: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_699, data_out=>output_MAC_2_699);
	MAC_2_700: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_700, data_out=>output_MAC_2_700);
	MAC_2_701: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_701, data_out=>output_MAC_2_701);
	MAC_2_702: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_702, data_out=>output_MAC_2_702);
	MAC_2_703: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_703, data_out=>output_MAC_2_703);
	MAC_2_704: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_704, data_out=>output_MAC_2_704);
	MAC_2_705: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_705, data_out=>output_MAC_2_705);
	MAC_2_706: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_706, data_out=>output_MAC_2_706);
	MAC_2_707: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_707, data_out=>output_MAC_2_707);
	MAC_2_708: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_708, data_out=>output_MAC_2_708);
	MAC_2_709: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_709, data_out=>output_MAC_2_709);
	MAC_2_710: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_710, data_out=>output_MAC_2_710);
	MAC_2_711: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_711, data_out=>output_MAC_2_711);
	MAC_2_712: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_712, data_out=>output_MAC_2_712);
	MAC_2_713: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_713, data_out=>output_MAC_2_713);
	MAC_2_714: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_714, data_out=>output_MAC_2_714);
	MAC_2_715: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_715, data_out=>output_MAC_2_715);
	MAC_2_716: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_716, data_out=>output_MAC_2_716);
	MAC_2_717: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_717, data_out=>output_MAC_2_717);
	MAC_2_718: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_718, data_out=>output_MAC_2_718);
	MAC_2_719: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_719, data_out=>output_MAC_2_719);
	MAC_2_720: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_720, data_out=>output_MAC_2_720);
	MAC_2_721: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_721, data_out=>output_MAC_2_721);
	MAC_2_722: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_722, data_out=>output_MAC_2_722);
	MAC_2_723: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_723, data_out=>output_MAC_2_723);
	MAC_2_724: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_724, data_out=>output_MAC_2_724);
	MAC_2_725: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_725, data_out=>output_MAC_2_725);
	MAC_2_726: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_726, data_out=>output_MAC_2_726);
	MAC_2_727: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_727, data_out=>output_MAC_2_727);
	MAC_2_728: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_728, data_out=>output_MAC_2_728);
	MAC_2_729: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_729, data_out=>output_MAC_2_729);
	MAC_2_730: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_730, data_out=>output_MAC_2_730);
	MAC_2_731: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_731, data_out=>output_MAC_2_731);
	MAC_2_732: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_732, data_out=>output_MAC_2_732);
	MAC_2_733: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_733, data_out=>output_MAC_2_733);
	MAC_2_734: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_734, data_out=>output_MAC_2_734);
	MAC_2_735: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_735, data_out=>output_MAC_2_735);
	MAC_2_736: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_736, data_out=>output_MAC_2_736);
	MAC_2_737: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_737, data_out=>output_MAC_2_737);
	MAC_2_738: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_738, data_out=>output_MAC_2_738);
	MAC_2_739: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_739, data_out=>output_MAC_2_739);
	MAC_2_740: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_740, data_out=>output_MAC_2_740);
	MAC_2_741: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_741, data_out=>output_MAC_2_741);
	MAC_2_742: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_742, data_out=>output_MAC_2_742);
	MAC_2_743: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_743, data_out=>output_MAC_2_743);
	MAC_2_744: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_744, data_out=>output_MAC_2_744);
	MAC_2_745: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_745, data_out=>output_MAC_2_745);
	MAC_2_746: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_746, data_out=>output_MAC_2_746);
	MAC_2_747: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_747, data_out=>output_MAC_2_747);
	MAC_2_748: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_748, data_out=>output_MAC_2_748);
	MAC_2_749: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_749, data_out=>output_MAC_2_749);
	MAC_2_750: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_750, data_out=>output_MAC_2_750);
	MAC_2_751: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_751, data_out=>output_MAC_2_751);
	MAC_2_752: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_752, data_out=>output_MAC_2_752);
	MAC_2_753: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_753, data_out=>output_MAC_2_753);
	MAC_2_754: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_754, data_out=>output_MAC_2_754);
	MAC_2_755: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_755, data_out=>output_MAC_2_755);
	MAC_2_756: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_756, data_out=>output_MAC_2_756);
	MAC_2_757: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_757, data_out=>output_MAC_2_757);
	MAC_2_758: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_758, data_out=>output_MAC_2_758);
	MAC_2_759: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_759, data_out=>output_MAC_2_759);
	MAC_2_760: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_760, data_out=>output_MAC_2_760);
	MAC_2_761: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_761, data_out=>output_MAC_2_761);
	MAC_2_762: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_762, data_out=>output_MAC_2_762);
	MAC_2_763: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_763, data_out=>output_MAC_2_763);
	MAC_2_764: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_764, data_out=>output_MAC_2_764);
	MAC_2_765: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_765, data_out=>output_MAC_2_765);
	MAC_2_766: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_766, data_out=>output_MAC_2_766);
	MAC_2_767: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_2, data_in_B=>input_col_767, data_out=>output_MAC_2_767);
	MAC_3_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_0, data_out=>output_MAC_3_0);
	MAC_3_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_1, data_out=>output_MAC_3_1);
	MAC_3_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_2, data_out=>output_MAC_3_2);
	MAC_3_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_3, data_out=>output_MAC_3_3);
	MAC_3_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_4, data_out=>output_MAC_3_4);
	MAC_3_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_5, data_out=>output_MAC_3_5);
	MAC_3_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_6, data_out=>output_MAC_3_6);
	MAC_3_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_7, data_out=>output_MAC_3_7);
	MAC_3_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_8, data_out=>output_MAC_3_8);
	MAC_3_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_9, data_out=>output_MAC_3_9);
	MAC_3_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_10, data_out=>output_MAC_3_10);
	MAC_3_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_11, data_out=>output_MAC_3_11);
	MAC_3_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_12, data_out=>output_MAC_3_12);
	MAC_3_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_13, data_out=>output_MAC_3_13);
	MAC_3_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_14, data_out=>output_MAC_3_14);
	MAC_3_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_15, data_out=>output_MAC_3_15);
	MAC_3_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_16, data_out=>output_MAC_3_16);
	MAC_3_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_17, data_out=>output_MAC_3_17);
	MAC_3_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_18, data_out=>output_MAC_3_18);
	MAC_3_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_19, data_out=>output_MAC_3_19);
	MAC_3_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_20, data_out=>output_MAC_3_20);
	MAC_3_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_21, data_out=>output_MAC_3_21);
	MAC_3_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_22, data_out=>output_MAC_3_22);
	MAC_3_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_23, data_out=>output_MAC_3_23);
	MAC_3_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_24, data_out=>output_MAC_3_24);
	MAC_3_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_25, data_out=>output_MAC_3_25);
	MAC_3_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_26, data_out=>output_MAC_3_26);
	MAC_3_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_27, data_out=>output_MAC_3_27);
	MAC_3_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_28, data_out=>output_MAC_3_28);
	MAC_3_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_29, data_out=>output_MAC_3_29);
	MAC_3_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_30, data_out=>output_MAC_3_30);
	MAC_3_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_31, data_out=>output_MAC_3_31);
	MAC_3_32: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_32, data_out=>output_MAC_3_32);
	MAC_3_33: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_33, data_out=>output_MAC_3_33);
	MAC_3_34: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_34, data_out=>output_MAC_3_34);
	MAC_3_35: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_35, data_out=>output_MAC_3_35);
	MAC_3_36: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_36, data_out=>output_MAC_3_36);
	MAC_3_37: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_37, data_out=>output_MAC_3_37);
	MAC_3_38: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_38, data_out=>output_MAC_3_38);
	MAC_3_39: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_39, data_out=>output_MAC_3_39);
	MAC_3_40: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_40, data_out=>output_MAC_3_40);
	MAC_3_41: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_41, data_out=>output_MAC_3_41);
	MAC_3_42: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_42, data_out=>output_MAC_3_42);
	MAC_3_43: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_43, data_out=>output_MAC_3_43);
	MAC_3_44: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_44, data_out=>output_MAC_3_44);
	MAC_3_45: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_45, data_out=>output_MAC_3_45);
	MAC_3_46: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_46, data_out=>output_MAC_3_46);
	MAC_3_47: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_47, data_out=>output_MAC_3_47);
	MAC_3_48: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_48, data_out=>output_MAC_3_48);
	MAC_3_49: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_49, data_out=>output_MAC_3_49);
	MAC_3_50: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_50, data_out=>output_MAC_3_50);
	MAC_3_51: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_51, data_out=>output_MAC_3_51);
	MAC_3_52: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_52, data_out=>output_MAC_3_52);
	MAC_3_53: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_53, data_out=>output_MAC_3_53);
	MAC_3_54: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_54, data_out=>output_MAC_3_54);
	MAC_3_55: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_55, data_out=>output_MAC_3_55);
	MAC_3_56: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_56, data_out=>output_MAC_3_56);
	MAC_3_57: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_57, data_out=>output_MAC_3_57);
	MAC_3_58: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_58, data_out=>output_MAC_3_58);
	MAC_3_59: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_59, data_out=>output_MAC_3_59);
	MAC_3_60: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_60, data_out=>output_MAC_3_60);
	MAC_3_61: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_61, data_out=>output_MAC_3_61);
	MAC_3_62: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_62, data_out=>output_MAC_3_62);
	MAC_3_63: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_63, data_out=>output_MAC_3_63);
	MAC_3_64: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_64, data_out=>output_MAC_3_64);
	MAC_3_65: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_65, data_out=>output_MAC_3_65);
	MAC_3_66: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_66, data_out=>output_MAC_3_66);
	MAC_3_67: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_67, data_out=>output_MAC_3_67);
	MAC_3_68: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_68, data_out=>output_MAC_3_68);
	MAC_3_69: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_69, data_out=>output_MAC_3_69);
	MAC_3_70: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_70, data_out=>output_MAC_3_70);
	MAC_3_71: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_71, data_out=>output_MAC_3_71);
	MAC_3_72: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_72, data_out=>output_MAC_3_72);
	MAC_3_73: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_73, data_out=>output_MAC_3_73);
	MAC_3_74: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_74, data_out=>output_MAC_3_74);
	MAC_3_75: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_75, data_out=>output_MAC_3_75);
	MAC_3_76: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_76, data_out=>output_MAC_3_76);
	MAC_3_77: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_77, data_out=>output_MAC_3_77);
	MAC_3_78: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_78, data_out=>output_MAC_3_78);
	MAC_3_79: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_79, data_out=>output_MAC_3_79);
	MAC_3_80: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_80, data_out=>output_MAC_3_80);
	MAC_3_81: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_81, data_out=>output_MAC_3_81);
	MAC_3_82: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_82, data_out=>output_MAC_3_82);
	MAC_3_83: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_83, data_out=>output_MAC_3_83);
	MAC_3_84: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_84, data_out=>output_MAC_3_84);
	MAC_3_85: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_85, data_out=>output_MAC_3_85);
	MAC_3_86: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_86, data_out=>output_MAC_3_86);
	MAC_3_87: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_87, data_out=>output_MAC_3_87);
	MAC_3_88: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_88, data_out=>output_MAC_3_88);
	MAC_3_89: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_89, data_out=>output_MAC_3_89);
	MAC_3_90: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_90, data_out=>output_MAC_3_90);
	MAC_3_91: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_91, data_out=>output_MAC_3_91);
	MAC_3_92: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_92, data_out=>output_MAC_3_92);
	MAC_3_93: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_93, data_out=>output_MAC_3_93);
	MAC_3_94: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_94, data_out=>output_MAC_3_94);
	MAC_3_95: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_95, data_out=>output_MAC_3_95);
	MAC_3_96: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_96, data_out=>output_MAC_3_96);
	MAC_3_97: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_97, data_out=>output_MAC_3_97);
	MAC_3_98: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_98, data_out=>output_MAC_3_98);
	MAC_3_99: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_99, data_out=>output_MAC_3_99);
	MAC_3_100: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_100, data_out=>output_MAC_3_100);
	MAC_3_101: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_101, data_out=>output_MAC_3_101);
	MAC_3_102: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_102, data_out=>output_MAC_3_102);
	MAC_3_103: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_103, data_out=>output_MAC_3_103);
	MAC_3_104: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_104, data_out=>output_MAC_3_104);
	MAC_3_105: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_105, data_out=>output_MAC_3_105);
	MAC_3_106: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_106, data_out=>output_MAC_3_106);
	MAC_3_107: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_107, data_out=>output_MAC_3_107);
	MAC_3_108: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_108, data_out=>output_MAC_3_108);
	MAC_3_109: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_109, data_out=>output_MAC_3_109);
	MAC_3_110: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_110, data_out=>output_MAC_3_110);
	MAC_3_111: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_111, data_out=>output_MAC_3_111);
	MAC_3_112: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_112, data_out=>output_MAC_3_112);
	MAC_3_113: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_113, data_out=>output_MAC_3_113);
	MAC_3_114: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_114, data_out=>output_MAC_3_114);
	MAC_3_115: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_115, data_out=>output_MAC_3_115);
	MAC_3_116: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_116, data_out=>output_MAC_3_116);
	MAC_3_117: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_117, data_out=>output_MAC_3_117);
	MAC_3_118: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_118, data_out=>output_MAC_3_118);
	MAC_3_119: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_119, data_out=>output_MAC_3_119);
	MAC_3_120: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_120, data_out=>output_MAC_3_120);
	MAC_3_121: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_121, data_out=>output_MAC_3_121);
	MAC_3_122: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_122, data_out=>output_MAC_3_122);
	MAC_3_123: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_123, data_out=>output_MAC_3_123);
	MAC_3_124: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_124, data_out=>output_MAC_3_124);
	MAC_3_125: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_125, data_out=>output_MAC_3_125);
	MAC_3_126: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_126, data_out=>output_MAC_3_126);
	MAC_3_127: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_127, data_out=>output_MAC_3_127);
	MAC_3_128: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_128, data_out=>output_MAC_3_128);
	MAC_3_129: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_129, data_out=>output_MAC_3_129);
	MAC_3_130: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_130, data_out=>output_MAC_3_130);
	MAC_3_131: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_131, data_out=>output_MAC_3_131);
	MAC_3_132: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_132, data_out=>output_MAC_3_132);
	MAC_3_133: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_133, data_out=>output_MAC_3_133);
	MAC_3_134: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_134, data_out=>output_MAC_3_134);
	MAC_3_135: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_135, data_out=>output_MAC_3_135);
	MAC_3_136: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_136, data_out=>output_MAC_3_136);
	MAC_3_137: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_137, data_out=>output_MAC_3_137);
	MAC_3_138: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_138, data_out=>output_MAC_3_138);
	MAC_3_139: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_139, data_out=>output_MAC_3_139);
	MAC_3_140: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_140, data_out=>output_MAC_3_140);
	MAC_3_141: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_141, data_out=>output_MAC_3_141);
	MAC_3_142: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_142, data_out=>output_MAC_3_142);
	MAC_3_143: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_143, data_out=>output_MAC_3_143);
	MAC_3_144: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_144, data_out=>output_MAC_3_144);
	MAC_3_145: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_145, data_out=>output_MAC_3_145);
	MAC_3_146: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_146, data_out=>output_MAC_3_146);
	MAC_3_147: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_147, data_out=>output_MAC_3_147);
	MAC_3_148: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_148, data_out=>output_MAC_3_148);
	MAC_3_149: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_149, data_out=>output_MAC_3_149);
	MAC_3_150: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_150, data_out=>output_MAC_3_150);
	MAC_3_151: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_151, data_out=>output_MAC_3_151);
	MAC_3_152: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_152, data_out=>output_MAC_3_152);
	MAC_3_153: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_153, data_out=>output_MAC_3_153);
	MAC_3_154: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_154, data_out=>output_MAC_3_154);
	MAC_3_155: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_155, data_out=>output_MAC_3_155);
	MAC_3_156: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_156, data_out=>output_MAC_3_156);
	MAC_3_157: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_157, data_out=>output_MAC_3_157);
	MAC_3_158: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_158, data_out=>output_MAC_3_158);
	MAC_3_159: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_159, data_out=>output_MAC_3_159);
	MAC_3_160: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_160, data_out=>output_MAC_3_160);
	MAC_3_161: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_161, data_out=>output_MAC_3_161);
	MAC_3_162: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_162, data_out=>output_MAC_3_162);
	MAC_3_163: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_163, data_out=>output_MAC_3_163);
	MAC_3_164: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_164, data_out=>output_MAC_3_164);
	MAC_3_165: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_165, data_out=>output_MAC_3_165);
	MAC_3_166: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_166, data_out=>output_MAC_3_166);
	MAC_3_167: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_167, data_out=>output_MAC_3_167);
	MAC_3_168: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_168, data_out=>output_MAC_3_168);
	MAC_3_169: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_169, data_out=>output_MAC_3_169);
	MAC_3_170: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_170, data_out=>output_MAC_3_170);
	MAC_3_171: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_171, data_out=>output_MAC_3_171);
	MAC_3_172: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_172, data_out=>output_MAC_3_172);
	MAC_3_173: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_173, data_out=>output_MAC_3_173);
	MAC_3_174: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_174, data_out=>output_MAC_3_174);
	MAC_3_175: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_175, data_out=>output_MAC_3_175);
	MAC_3_176: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_176, data_out=>output_MAC_3_176);
	MAC_3_177: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_177, data_out=>output_MAC_3_177);
	MAC_3_178: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_178, data_out=>output_MAC_3_178);
	MAC_3_179: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_179, data_out=>output_MAC_3_179);
	MAC_3_180: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_180, data_out=>output_MAC_3_180);
	MAC_3_181: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_181, data_out=>output_MAC_3_181);
	MAC_3_182: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_182, data_out=>output_MAC_3_182);
	MAC_3_183: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_183, data_out=>output_MAC_3_183);
	MAC_3_184: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_184, data_out=>output_MAC_3_184);
	MAC_3_185: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_185, data_out=>output_MAC_3_185);
	MAC_3_186: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_186, data_out=>output_MAC_3_186);
	MAC_3_187: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_187, data_out=>output_MAC_3_187);
	MAC_3_188: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_188, data_out=>output_MAC_3_188);
	MAC_3_189: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_189, data_out=>output_MAC_3_189);
	MAC_3_190: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_190, data_out=>output_MAC_3_190);
	MAC_3_191: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_191, data_out=>output_MAC_3_191);
	MAC_3_192: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_192, data_out=>output_MAC_3_192);
	MAC_3_193: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_193, data_out=>output_MAC_3_193);
	MAC_3_194: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_194, data_out=>output_MAC_3_194);
	MAC_3_195: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_195, data_out=>output_MAC_3_195);
	MAC_3_196: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_196, data_out=>output_MAC_3_196);
	MAC_3_197: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_197, data_out=>output_MAC_3_197);
	MAC_3_198: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_198, data_out=>output_MAC_3_198);
	MAC_3_199: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_199, data_out=>output_MAC_3_199);
	MAC_3_200: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_200, data_out=>output_MAC_3_200);
	MAC_3_201: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_201, data_out=>output_MAC_3_201);
	MAC_3_202: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_202, data_out=>output_MAC_3_202);
	MAC_3_203: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_203, data_out=>output_MAC_3_203);
	MAC_3_204: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_204, data_out=>output_MAC_3_204);
	MAC_3_205: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_205, data_out=>output_MAC_3_205);
	MAC_3_206: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_206, data_out=>output_MAC_3_206);
	MAC_3_207: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_207, data_out=>output_MAC_3_207);
	MAC_3_208: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_208, data_out=>output_MAC_3_208);
	MAC_3_209: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_209, data_out=>output_MAC_3_209);
	MAC_3_210: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_210, data_out=>output_MAC_3_210);
	MAC_3_211: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_211, data_out=>output_MAC_3_211);
	MAC_3_212: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_212, data_out=>output_MAC_3_212);
	MAC_3_213: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_213, data_out=>output_MAC_3_213);
	MAC_3_214: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_214, data_out=>output_MAC_3_214);
	MAC_3_215: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_215, data_out=>output_MAC_3_215);
	MAC_3_216: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_216, data_out=>output_MAC_3_216);
	MAC_3_217: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_217, data_out=>output_MAC_3_217);
	MAC_3_218: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_218, data_out=>output_MAC_3_218);
	MAC_3_219: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_219, data_out=>output_MAC_3_219);
	MAC_3_220: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_220, data_out=>output_MAC_3_220);
	MAC_3_221: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_221, data_out=>output_MAC_3_221);
	MAC_3_222: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_222, data_out=>output_MAC_3_222);
	MAC_3_223: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_223, data_out=>output_MAC_3_223);
	MAC_3_224: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_224, data_out=>output_MAC_3_224);
	MAC_3_225: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_225, data_out=>output_MAC_3_225);
	MAC_3_226: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_226, data_out=>output_MAC_3_226);
	MAC_3_227: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_227, data_out=>output_MAC_3_227);
	MAC_3_228: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_228, data_out=>output_MAC_3_228);
	MAC_3_229: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_229, data_out=>output_MAC_3_229);
	MAC_3_230: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_230, data_out=>output_MAC_3_230);
	MAC_3_231: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_231, data_out=>output_MAC_3_231);
	MAC_3_232: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_232, data_out=>output_MAC_3_232);
	MAC_3_233: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_233, data_out=>output_MAC_3_233);
	MAC_3_234: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_234, data_out=>output_MAC_3_234);
	MAC_3_235: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_235, data_out=>output_MAC_3_235);
	MAC_3_236: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_236, data_out=>output_MAC_3_236);
	MAC_3_237: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_237, data_out=>output_MAC_3_237);
	MAC_3_238: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_238, data_out=>output_MAC_3_238);
	MAC_3_239: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_239, data_out=>output_MAC_3_239);
	MAC_3_240: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_240, data_out=>output_MAC_3_240);
	MAC_3_241: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_241, data_out=>output_MAC_3_241);
	MAC_3_242: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_242, data_out=>output_MAC_3_242);
	MAC_3_243: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_243, data_out=>output_MAC_3_243);
	MAC_3_244: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_244, data_out=>output_MAC_3_244);
	MAC_3_245: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_245, data_out=>output_MAC_3_245);
	MAC_3_246: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_246, data_out=>output_MAC_3_246);
	MAC_3_247: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_247, data_out=>output_MAC_3_247);
	MAC_3_248: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_248, data_out=>output_MAC_3_248);
	MAC_3_249: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_249, data_out=>output_MAC_3_249);
	MAC_3_250: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_250, data_out=>output_MAC_3_250);
	MAC_3_251: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_251, data_out=>output_MAC_3_251);
	MAC_3_252: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_252, data_out=>output_MAC_3_252);
	MAC_3_253: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_253, data_out=>output_MAC_3_253);
	MAC_3_254: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_254, data_out=>output_MAC_3_254);
	MAC_3_255: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_255, data_out=>output_MAC_3_255);
	MAC_3_256: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_256, data_out=>output_MAC_3_256);
	MAC_3_257: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_257, data_out=>output_MAC_3_257);
	MAC_3_258: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_258, data_out=>output_MAC_3_258);
	MAC_3_259: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_259, data_out=>output_MAC_3_259);
	MAC_3_260: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_260, data_out=>output_MAC_3_260);
	MAC_3_261: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_261, data_out=>output_MAC_3_261);
	MAC_3_262: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_262, data_out=>output_MAC_3_262);
	MAC_3_263: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_263, data_out=>output_MAC_3_263);
	MAC_3_264: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_264, data_out=>output_MAC_3_264);
	MAC_3_265: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_265, data_out=>output_MAC_3_265);
	MAC_3_266: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_266, data_out=>output_MAC_3_266);
	MAC_3_267: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_267, data_out=>output_MAC_3_267);
	MAC_3_268: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_268, data_out=>output_MAC_3_268);
	MAC_3_269: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_269, data_out=>output_MAC_3_269);
	MAC_3_270: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_270, data_out=>output_MAC_3_270);
	MAC_3_271: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_271, data_out=>output_MAC_3_271);
	MAC_3_272: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_272, data_out=>output_MAC_3_272);
	MAC_3_273: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_273, data_out=>output_MAC_3_273);
	MAC_3_274: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_274, data_out=>output_MAC_3_274);
	MAC_3_275: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_275, data_out=>output_MAC_3_275);
	MAC_3_276: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_276, data_out=>output_MAC_3_276);
	MAC_3_277: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_277, data_out=>output_MAC_3_277);
	MAC_3_278: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_278, data_out=>output_MAC_3_278);
	MAC_3_279: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_279, data_out=>output_MAC_3_279);
	MAC_3_280: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_280, data_out=>output_MAC_3_280);
	MAC_3_281: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_281, data_out=>output_MAC_3_281);
	MAC_3_282: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_282, data_out=>output_MAC_3_282);
	MAC_3_283: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_283, data_out=>output_MAC_3_283);
	MAC_3_284: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_284, data_out=>output_MAC_3_284);
	MAC_3_285: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_285, data_out=>output_MAC_3_285);
	MAC_3_286: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_286, data_out=>output_MAC_3_286);
	MAC_3_287: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_287, data_out=>output_MAC_3_287);
	MAC_3_288: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_288, data_out=>output_MAC_3_288);
	MAC_3_289: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_289, data_out=>output_MAC_3_289);
	MAC_3_290: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_290, data_out=>output_MAC_3_290);
	MAC_3_291: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_291, data_out=>output_MAC_3_291);
	MAC_3_292: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_292, data_out=>output_MAC_3_292);
	MAC_3_293: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_293, data_out=>output_MAC_3_293);
	MAC_3_294: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_294, data_out=>output_MAC_3_294);
	MAC_3_295: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_295, data_out=>output_MAC_3_295);
	MAC_3_296: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_296, data_out=>output_MAC_3_296);
	MAC_3_297: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_297, data_out=>output_MAC_3_297);
	MAC_3_298: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_298, data_out=>output_MAC_3_298);
	MAC_3_299: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_299, data_out=>output_MAC_3_299);
	MAC_3_300: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_300, data_out=>output_MAC_3_300);
	MAC_3_301: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_301, data_out=>output_MAC_3_301);
	MAC_3_302: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_302, data_out=>output_MAC_3_302);
	MAC_3_303: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_303, data_out=>output_MAC_3_303);
	MAC_3_304: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_304, data_out=>output_MAC_3_304);
	MAC_3_305: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_305, data_out=>output_MAC_3_305);
	MAC_3_306: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_306, data_out=>output_MAC_3_306);
	MAC_3_307: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_307, data_out=>output_MAC_3_307);
	MAC_3_308: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_308, data_out=>output_MAC_3_308);
	MAC_3_309: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_309, data_out=>output_MAC_3_309);
	MAC_3_310: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_310, data_out=>output_MAC_3_310);
	MAC_3_311: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_311, data_out=>output_MAC_3_311);
	MAC_3_312: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_312, data_out=>output_MAC_3_312);
	MAC_3_313: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_313, data_out=>output_MAC_3_313);
	MAC_3_314: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_314, data_out=>output_MAC_3_314);
	MAC_3_315: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_315, data_out=>output_MAC_3_315);
	MAC_3_316: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_316, data_out=>output_MAC_3_316);
	MAC_3_317: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_317, data_out=>output_MAC_3_317);
	MAC_3_318: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_318, data_out=>output_MAC_3_318);
	MAC_3_319: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_319, data_out=>output_MAC_3_319);
	MAC_3_320: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_320, data_out=>output_MAC_3_320);
	MAC_3_321: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_321, data_out=>output_MAC_3_321);
	MAC_3_322: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_322, data_out=>output_MAC_3_322);
	MAC_3_323: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_323, data_out=>output_MAC_3_323);
	MAC_3_324: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_324, data_out=>output_MAC_3_324);
	MAC_3_325: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_325, data_out=>output_MAC_3_325);
	MAC_3_326: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_326, data_out=>output_MAC_3_326);
	MAC_3_327: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_327, data_out=>output_MAC_3_327);
	MAC_3_328: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_328, data_out=>output_MAC_3_328);
	MAC_3_329: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_329, data_out=>output_MAC_3_329);
	MAC_3_330: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_330, data_out=>output_MAC_3_330);
	MAC_3_331: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_331, data_out=>output_MAC_3_331);
	MAC_3_332: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_332, data_out=>output_MAC_3_332);
	MAC_3_333: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_333, data_out=>output_MAC_3_333);
	MAC_3_334: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_334, data_out=>output_MAC_3_334);
	MAC_3_335: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_335, data_out=>output_MAC_3_335);
	MAC_3_336: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_336, data_out=>output_MAC_3_336);
	MAC_3_337: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_337, data_out=>output_MAC_3_337);
	MAC_3_338: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_338, data_out=>output_MAC_3_338);
	MAC_3_339: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_339, data_out=>output_MAC_3_339);
	MAC_3_340: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_340, data_out=>output_MAC_3_340);
	MAC_3_341: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_341, data_out=>output_MAC_3_341);
	MAC_3_342: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_342, data_out=>output_MAC_3_342);
	MAC_3_343: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_343, data_out=>output_MAC_3_343);
	MAC_3_344: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_344, data_out=>output_MAC_3_344);
	MAC_3_345: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_345, data_out=>output_MAC_3_345);
	MAC_3_346: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_346, data_out=>output_MAC_3_346);
	MAC_3_347: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_347, data_out=>output_MAC_3_347);
	MAC_3_348: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_348, data_out=>output_MAC_3_348);
	MAC_3_349: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_349, data_out=>output_MAC_3_349);
	MAC_3_350: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_350, data_out=>output_MAC_3_350);
	MAC_3_351: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_351, data_out=>output_MAC_3_351);
	MAC_3_352: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_352, data_out=>output_MAC_3_352);
	MAC_3_353: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_353, data_out=>output_MAC_3_353);
	MAC_3_354: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_354, data_out=>output_MAC_3_354);
	MAC_3_355: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_355, data_out=>output_MAC_3_355);
	MAC_3_356: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_356, data_out=>output_MAC_3_356);
	MAC_3_357: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_357, data_out=>output_MAC_3_357);
	MAC_3_358: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_358, data_out=>output_MAC_3_358);
	MAC_3_359: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_359, data_out=>output_MAC_3_359);
	MAC_3_360: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_360, data_out=>output_MAC_3_360);
	MAC_3_361: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_361, data_out=>output_MAC_3_361);
	MAC_3_362: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_362, data_out=>output_MAC_3_362);
	MAC_3_363: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_363, data_out=>output_MAC_3_363);
	MAC_3_364: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_364, data_out=>output_MAC_3_364);
	MAC_3_365: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_365, data_out=>output_MAC_3_365);
	MAC_3_366: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_366, data_out=>output_MAC_3_366);
	MAC_3_367: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_367, data_out=>output_MAC_3_367);
	MAC_3_368: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_368, data_out=>output_MAC_3_368);
	MAC_3_369: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_369, data_out=>output_MAC_3_369);
	MAC_3_370: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_370, data_out=>output_MAC_3_370);
	MAC_3_371: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_371, data_out=>output_MAC_3_371);
	MAC_3_372: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_372, data_out=>output_MAC_3_372);
	MAC_3_373: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_373, data_out=>output_MAC_3_373);
	MAC_3_374: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_374, data_out=>output_MAC_3_374);
	MAC_3_375: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_375, data_out=>output_MAC_3_375);
	MAC_3_376: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_376, data_out=>output_MAC_3_376);
	MAC_3_377: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_377, data_out=>output_MAC_3_377);
	MAC_3_378: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_378, data_out=>output_MAC_3_378);
	MAC_3_379: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_379, data_out=>output_MAC_3_379);
	MAC_3_380: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_380, data_out=>output_MAC_3_380);
	MAC_3_381: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_381, data_out=>output_MAC_3_381);
	MAC_3_382: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_382, data_out=>output_MAC_3_382);
	MAC_3_383: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_383, data_out=>output_MAC_3_383);
	MAC_3_384: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_384, data_out=>output_MAC_3_384);
	MAC_3_385: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_385, data_out=>output_MAC_3_385);
	MAC_3_386: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_386, data_out=>output_MAC_3_386);
	MAC_3_387: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_387, data_out=>output_MAC_3_387);
	MAC_3_388: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_388, data_out=>output_MAC_3_388);
	MAC_3_389: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_389, data_out=>output_MAC_3_389);
	MAC_3_390: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_390, data_out=>output_MAC_3_390);
	MAC_3_391: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_391, data_out=>output_MAC_3_391);
	MAC_3_392: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_392, data_out=>output_MAC_3_392);
	MAC_3_393: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_393, data_out=>output_MAC_3_393);
	MAC_3_394: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_394, data_out=>output_MAC_3_394);
	MAC_3_395: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_395, data_out=>output_MAC_3_395);
	MAC_3_396: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_396, data_out=>output_MAC_3_396);
	MAC_3_397: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_397, data_out=>output_MAC_3_397);
	MAC_3_398: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_398, data_out=>output_MAC_3_398);
	MAC_3_399: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_399, data_out=>output_MAC_3_399);
	MAC_3_400: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_400, data_out=>output_MAC_3_400);
	MAC_3_401: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_401, data_out=>output_MAC_3_401);
	MAC_3_402: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_402, data_out=>output_MAC_3_402);
	MAC_3_403: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_403, data_out=>output_MAC_3_403);
	MAC_3_404: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_404, data_out=>output_MAC_3_404);
	MAC_3_405: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_405, data_out=>output_MAC_3_405);
	MAC_3_406: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_406, data_out=>output_MAC_3_406);
	MAC_3_407: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_407, data_out=>output_MAC_3_407);
	MAC_3_408: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_408, data_out=>output_MAC_3_408);
	MAC_3_409: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_409, data_out=>output_MAC_3_409);
	MAC_3_410: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_410, data_out=>output_MAC_3_410);
	MAC_3_411: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_411, data_out=>output_MAC_3_411);
	MAC_3_412: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_412, data_out=>output_MAC_3_412);
	MAC_3_413: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_413, data_out=>output_MAC_3_413);
	MAC_3_414: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_414, data_out=>output_MAC_3_414);
	MAC_3_415: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_415, data_out=>output_MAC_3_415);
	MAC_3_416: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_416, data_out=>output_MAC_3_416);
	MAC_3_417: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_417, data_out=>output_MAC_3_417);
	MAC_3_418: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_418, data_out=>output_MAC_3_418);
	MAC_3_419: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_419, data_out=>output_MAC_3_419);
	MAC_3_420: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_420, data_out=>output_MAC_3_420);
	MAC_3_421: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_421, data_out=>output_MAC_3_421);
	MAC_3_422: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_422, data_out=>output_MAC_3_422);
	MAC_3_423: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_423, data_out=>output_MAC_3_423);
	MAC_3_424: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_424, data_out=>output_MAC_3_424);
	MAC_3_425: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_425, data_out=>output_MAC_3_425);
	MAC_3_426: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_426, data_out=>output_MAC_3_426);
	MAC_3_427: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_427, data_out=>output_MAC_3_427);
	MAC_3_428: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_428, data_out=>output_MAC_3_428);
	MAC_3_429: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_429, data_out=>output_MAC_3_429);
	MAC_3_430: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_430, data_out=>output_MAC_3_430);
	MAC_3_431: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_431, data_out=>output_MAC_3_431);
	MAC_3_432: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_432, data_out=>output_MAC_3_432);
	MAC_3_433: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_433, data_out=>output_MAC_3_433);
	MAC_3_434: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_434, data_out=>output_MAC_3_434);
	MAC_3_435: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_435, data_out=>output_MAC_3_435);
	MAC_3_436: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_436, data_out=>output_MAC_3_436);
	MAC_3_437: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_437, data_out=>output_MAC_3_437);
	MAC_3_438: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_438, data_out=>output_MAC_3_438);
	MAC_3_439: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_439, data_out=>output_MAC_3_439);
	MAC_3_440: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_440, data_out=>output_MAC_3_440);
	MAC_3_441: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_441, data_out=>output_MAC_3_441);
	MAC_3_442: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_442, data_out=>output_MAC_3_442);
	MAC_3_443: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_443, data_out=>output_MAC_3_443);
	MAC_3_444: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_444, data_out=>output_MAC_3_444);
	MAC_3_445: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_445, data_out=>output_MAC_3_445);
	MAC_3_446: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_446, data_out=>output_MAC_3_446);
	MAC_3_447: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_447, data_out=>output_MAC_3_447);
	MAC_3_448: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_448, data_out=>output_MAC_3_448);
	MAC_3_449: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_449, data_out=>output_MAC_3_449);
	MAC_3_450: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_450, data_out=>output_MAC_3_450);
	MAC_3_451: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_451, data_out=>output_MAC_3_451);
	MAC_3_452: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_452, data_out=>output_MAC_3_452);
	MAC_3_453: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_453, data_out=>output_MAC_3_453);
	MAC_3_454: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_454, data_out=>output_MAC_3_454);
	MAC_3_455: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_455, data_out=>output_MAC_3_455);
	MAC_3_456: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_456, data_out=>output_MAC_3_456);
	MAC_3_457: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_457, data_out=>output_MAC_3_457);
	MAC_3_458: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_458, data_out=>output_MAC_3_458);
	MAC_3_459: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_459, data_out=>output_MAC_3_459);
	MAC_3_460: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_460, data_out=>output_MAC_3_460);
	MAC_3_461: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_461, data_out=>output_MAC_3_461);
	MAC_3_462: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_462, data_out=>output_MAC_3_462);
	MAC_3_463: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_463, data_out=>output_MAC_3_463);
	MAC_3_464: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_464, data_out=>output_MAC_3_464);
	MAC_3_465: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_465, data_out=>output_MAC_3_465);
	MAC_3_466: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_466, data_out=>output_MAC_3_466);
	MAC_3_467: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_467, data_out=>output_MAC_3_467);
	MAC_3_468: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_468, data_out=>output_MAC_3_468);
	MAC_3_469: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_469, data_out=>output_MAC_3_469);
	MAC_3_470: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_470, data_out=>output_MAC_3_470);
	MAC_3_471: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_471, data_out=>output_MAC_3_471);
	MAC_3_472: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_472, data_out=>output_MAC_3_472);
	MAC_3_473: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_473, data_out=>output_MAC_3_473);
	MAC_3_474: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_474, data_out=>output_MAC_3_474);
	MAC_3_475: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_475, data_out=>output_MAC_3_475);
	MAC_3_476: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_476, data_out=>output_MAC_3_476);
	MAC_3_477: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_477, data_out=>output_MAC_3_477);
	MAC_3_478: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_478, data_out=>output_MAC_3_478);
	MAC_3_479: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_479, data_out=>output_MAC_3_479);
	MAC_3_480: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_480, data_out=>output_MAC_3_480);
	MAC_3_481: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_481, data_out=>output_MAC_3_481);
	MAC_3_482: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_482, data_out=>output_MAC_3_482);
	MAC_3_483: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_483, data_out=>output_MAC_3_483);
	MAC_3_484: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_484, data_out=>output_MAC_3_484);
	MAC_3_485: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_485, data_out=>output_MAC_3_485);
	MAC_3_486: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_486, data_out=>output_MAC_3_486);
	MAC_3_487: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_487, data_out=>output_MAC_3_487);
	MAC_3_488: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_488, data_out=>output_MAC_3_488);
	MAC_3_489: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_489, data_out=>output_MAC_3_489);
	MAC_3_490: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_490, data_out=>output_MAC_3_490);
	MAC_3_491: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_491, data_out=>output_MAC_3_491);
	MAC_3_492: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_492, data_out=>output_MAC_3_492);
	MAC_3_493: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_493, data_out=>output_MAC_3_493);
	MAC_3_494: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_494, data_out=>output_MAC_3_494);
	MAC_3_495: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_495, data_out=>output_MAC_3_495);
	MAC_3_496: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_496, data_out=>output_MAC_3_496);
	MAC_3_497: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_497, data_out=>output_MAC_3_497);
	MAC_3_498: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_498, data_out=>output_MAC_3_498);
	MAC_3_499: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_499, data_out=>output_MAC_3_499);
	MAC_3_500: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_500, data_out=>output_MAC_3_500);
	MAC_3_501: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_501, data_out=>output_MAC_3_501);
	MAC_3_502: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_502, data_out=>output_MAC_3_502);
	MAC_3_503: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_503, data_out=>output_MAC_3_503);
	MAC_3_504: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_504, data_out=>output_MAC_3_504);
	MAC_3_505: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_505, data_out=>output_MAC_3_505);
	MAC_3_506: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_506, data_out=>output_MAC_3_506);
	MAC_3_507: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_507, data_out=>output_MAC_3_507);
	MAC_3_508: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_508, data_out=>output_MAC_3_508);
	MAC_3_509: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_509, data_out=>output_MAC_3_509);
	MAC_3_510: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_510, data_out=>output_MAC_3_510);
	MAC_3_511: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_511, data_out=>output_MAC_3_511);
	MAC_3_512: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_512, data_out=>output_MAC_3_512);
	MAC_3_513: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_513, data_out=>output_MAC_3_513);
	MAC_3_514: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_514, data_out=>output_MAC_3_514);
	MAC_3_515: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_515, data_out=>output_MAC_3_515);
	MAC_3_516: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_516, data_out=>output_MAC_3_516);
	MAC_3_517: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_517, data_out=>output_MAC_3_517);
	MAC_3_518: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_518, data_out=>output_MAC_3_518);
	MAC_3_519: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_519, data_out=>output_MAC_3_519);
	MAC_3_520: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_520, data_out=>output_MAC_3_520);
	MAC_3_521: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_521, data_out=>output_MAC_3_521);
	MAC_3_522: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_522, data_out=>output_MAC_3_522);
	MAC_3_523: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_523, data_out=>output_MAC_3_523);
	MAC_3_524: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_524, data_out=>output_MAC_3_524);
	MAC_3_525: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_525, data_out=>output_MAC_3_525);
	MAC_3_526: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_526, data_out=>output_MAC_3_526);
	MAC_3_527: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_527, data_out=>output_MAC_3_527);
	MAC_3_528: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_528, data_out=>output_MAC_3_528);
	MAC_3_529: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_529, data_out=>output_MAC_3_529);
	MAC_3_530: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_530, data_out=>output_MAC_3_530);
	MAC_3_531: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_531, data_out=>output_MAC_3_531);
	MAC_3_532: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_532, data_out=>output_MAC_3_532);
	MAC_3_533: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_533, data_out=>output_MAC_3_533);
	MAC_3_534: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_534, data_out=>output_MAC_3_534);
	MAC_3_535: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_535, data_out=>output_MAC_3_535);
	MAC_3_536: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_536, data_out=>output_MAC_3_536);
	MAC_3_537: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_537, data_out=>output_MAC_3_537);
	MAC_3_538: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_538, data_out=>output_MAC_3_538);
	MAC_3_539: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_539, data_out=>output_MAC_3_539);
	MAC_3_540: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_540, data_out=>output_MAC_3_540);
	MAC_3_541: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_541, data_out=>output_MAC_3_541);
	MAC_3_542: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_542, data_out=>output_MAC_3_542);
	MAC_3_543: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_543, data_out=>output_MAC_3_543);
	MAC_3_544: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_544, data_out=>output_MAC_3_544);
	MAC_3_545: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_545, data_out=>output_MAC_3_545);
	MAC_3_546: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_546, data_out=>output_MAC_3_546);
	MAC_3_547: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_547, data_out=>output_MAC_3_547);
	MAC_3_548: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_548, data_out=>output_MAC_3_548);
	MAC_3_549: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_549, data_out=>output_MAC_3_549);
	MAC_3_550: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_550, data_out=>output_MAC_3_550);
	MAC_3_551: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_551, data_out=>output_MAC_3_551);
	MAC_3_552: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_552, data_out=>output_MAC_3_552);
	MAC_3_553: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_553, data_out=>output_MAC_3_553);
	MAC_3_554: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_554, data_out=>output_MAC_3_554);
	MAC_3_555: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_555, data_out=>output_MAC_3_555);
	MAC_3_556: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_556, data_out=>output_MAC_3_556);
	MAC_3_557: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_557, data_out=>output_MAC_3_557);
	MAC_3_558: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_558, data_out=>output_MAC_3_558);
	MAC_3_559: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_559, data_out=>output_MAC_3_559);
	MAC_3_560: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_560, data_out=>output_MAC_3_560);
	MAC_3_561: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_561, data_out=>output_MAC_3_561);
	MAC_3_562: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_562, data_out=>output_MAC_3_562);
	MAC_3_563: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_563, data_out=>output_MAC_3_563);
	MAC_3_564: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_564, data_out=>output_MAC_3_564);
	MAC_3_565: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_565, data_out=>output_MAC_3_565);
	MAC_3_566: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_566, data_out=>output_MAC_3_566);
	MAC_3_567: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_567, data_out=>output_MAC_3_567);
	MAC_3_568: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_568, data_out=>output_MAC_3_568);
	MAC_3_569: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_569, data_out=>output_MAC_3_569);
	MAC_3_570: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_570, data_out=>output_MAC_3_570);
	MAC_3_571: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_571, data_out=>output_MAC_3_571);
	MAC_3_572: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_572, data_out=>output_MAC_3_572);
	MAC_3_573: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_573, data_out=>output_MAC_3_573);
	MAC_3_574: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_574, data_out=>output_MAC_3_574);
	MAC_3_575: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_575, data_out=>output_MAC_3_575);
	MAC_3_576: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_576, data_out=>output_MAC_3_576);
	MAC_3_577: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_577, data_out=>output_MAC_3_577);
	MAC_3_578: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_578, data_out=>output_MAC_3_578);
	MAC_3_579: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_579, data_out=>output_MAC_3_579);
	MAC_3_580: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_580, data_out=>output_MAC_3_580);
	MAC_3_581: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_581, data_out=>output_MAC_3_581);
	MAC_3_582: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_582, data_out=>output_MAC_3_582);
	MAC_3_583: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_583, data_out=>output_MAC_3_583);
	MAC_3_584: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_584, data_out=>output_MAC_3_584);
	MAC_3_585: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_585, data_out=>output_MAC_3_585);
	MAC_3_586: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_586, data_out=>output_MAC_3_586);
	MAC_3_587: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_587, data_out=>output_MAC_3_587);
	MAC_3_588: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_588, data_out=>output_MAC_3_588);
	MAC_3_589: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_589, data_out=>output_MAC_3_589);
	MAC_3_590: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_590, data_out=>output_MAC_3_590);
	MAC_3_591: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_591, data_out=>output_MAC_3_591);
	MAC_3_592: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_592, data_out=>output_MAC_3_592);
	MAC_3_593: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_593, data_out=>output_MAC_3_593);
	MAC_3_594: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_594, data_out=>output_MAC_3_594);
	MAC_3_595: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_595, data_out=>output_MAC_3_595);
	MAC_3_596: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_596, data_out=>output_MAC_3_596);
	MAC_3_597: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_597, data_out=>output_MAC_3_597);
	MAC_3_598: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_598, data_out=>output_MAC_3_598);
	MAC_3_599: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_599, data_out=>output_MAC_3_599);
	MAC_3_600: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_600, data_out=>output_MAC_3_600);
	MAC_3_601: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_601, data_out=>output_MAC_3_601);
	MAC_3_602: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_602, data_out=>output_MAC_3_602);
	MAC_3_603: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_603, data_out=>output_MAC_3_603);
	MAC_3_604: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_604, data_out=>output_MAC_3_604);
	MAC_3_605: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_605, data_out=>output_MAC_3_605);
	MAC_3_606: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_606, data_out=>output_MAC_3_606);
	MAC_3_607: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_607, data_out=>output_MAC_3_607);
	MAC_3_608: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_608, data_out=>output_MAC_3_608);
	MAC_3_609: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_609, data_out=>output_MAC_3_609);
	MAC_3_610: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_610, data_out=>output_MAC_3_610);
	MAC_3_611: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_611, data_out=>output_MAC_3_611);
	MAC_3_612: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_612, data_out=>output_MAC_3_612);
	MAC_3_613: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_613, data_out=>output_MAC_3_613);
	MAC_3_614: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_614, data_out=>output_MAC_3_614);
	MAC_3_615: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_615, data_out=>output_MAC_3_615);
	MAC_3_616: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_616, data_out=>output_MAC_3_616);
	MAC_3_617: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_617, data_out=>output_MAC_3_617);
	MAC_3_618: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_618, data_out=>output_MAC_3_618);
	MAC_3_619: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_619, data_out=>output_MAC_3_619);
	MAC_3_620: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_620, data_out=>output_MAC_3_620);
	MAC_3_621: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_621, data_out=>output_MAC_3_621);
	MAC_3_622: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_622, data_out=>output_MAC_3_622);
	MAC_3_623: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_623, data_out=>output_MAC_3_623);
	MAC_3_624: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_624, data_out=>output_MAC_3_624);
	MAC_3_625: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_625, data_out=>output_MAC_3_625);
	MAC_3_626: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_626, data_out=>output_MAC_3_626);
	MAC_3_627: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_627, data_out=>output_MAC_3_627);
	MAC_3_628: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_628, data_out=>output_MAC_3_628);
	MAC_3_629: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_629, data_out=>output_MAC_3_629);
	MAC_3_630: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_630, data_out=>output_MAC_3_630);
	MAC_3_631: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_631, data_out=>output_MAC_3_631);
	MAC_3_632: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_632, data_out=>output_MAC_3_632);
	MAC_3_633: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_633, data_out=>output_MAC_3_633);
	MAC_3_634: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_634, data_out=>output_MAC_3_634);
	MAC_3_635: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_635, data_out=>output_MAC_3_635);
	MAC_3_636: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_636, data_out=>output_MAC_3_636);
	MAC_3_637: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_637, data_out=>output_MAC_3_637);
	MAC_3_638: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_638, data_out=>output_MAC_3_638);
	MAC_3_639: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_639, data_out=>output_MAC_3_639);
	MAC_3_640: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_640, data_out=>output_MAC_3_640);
	MAC_3_641: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_641, data_out=>output_MAC_3_641);
	MAC_3_642: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_642, data_out=>output_MAC_3_642);
	MAC_3_643: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_643, data_out=>output_MAC_3_643);
	MAC_3_644: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_644, data_out=>output_MAC_3_644);
	MAC_3_645: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_645, data_out=>output_MAC_3_645);
	MAC_3_646: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_646, data_out=>output_MAC_3_646);
	MAC_3_647: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_647, data_out=>output_MAC_3_647);
	MAC_3_648: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_648, data_out=>output_MAC_3_648);
	MAC_3_649: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_649, data_out=>output_MAC_3_649);
	MAC_3_650: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_650, data_out=>output_MAC_3_650);
	MAC_3_651: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_651, data_out=>output_MAC_3_651);
	MAC_3_652: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_652, data_out=>output_MAC_3_652);
	MAC_3_653: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_653, data_out=>output_MAC_3_653);
	MAC_3_654: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_654, data_out=>output_MAC_3_654);
	MAC_3_655: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_655, data_out=>output_MAC_3_655);
	MAC_3_656: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_656, data_out=>output_MAC_3_656);
	MAC_3_657: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_657, data_out=>output_MAC_3_657);
	MAC_3_658: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_658, data_out=>output_MAC_3_658);
	MAC_3_659: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_659, data_out=>output_MAC_3_659);
	MAC_3_660: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_660, data_out=>output_MAC_3_660);
	MAC_3_661: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_661, data_out=>output_MAC_3_661);
	MAC_3_662: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_662, data_out=>output_MAC_3_662);
	MAC_3_663: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_663, data_out=>output_MAC_3_663);
	MAC_3_664: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_664, data_out=>output_MAC_3_664);
	MAC_3_665: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_665, data_out=>output_MAC_3_665);
	MAC_3_666: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_666, data_out=>output_MAC_3_666);
	MAC_3_667: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_667, data_out=>output_MAC_3_667);
	MAC_3_668: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_668, data_out=>output_MAC_3_668);
	MAC_3_669: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_669, data_out=>output_MAC_3_669);
	MAC_3_670: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_670, data_out=>output_MAC_3_670);
	MAC_3_671: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_671, data_out=>output_MAC_3_671);
	MAC_3_672: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_672, data_out=>output_MAC_3_672);
	MAC_3_673: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_673, data_out=>output_MAC_3_673);
	MAC_3_674: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_674, data_out=>output_MAC_3_674);
	MAC_3_675: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_675, data_out=>output_MAC_3_675);
	MAC_3_676: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_676, data_out=>output_MAC_3_676);
	MAC_3_677: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_677, data_out=>output_MAC_3_677);
	MAC_3_678: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_678, data_out=>output_MAC_3_678);
	MAC_3_679: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_679, data_out=>output_MAC_3_679);
	MAC_3_680: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_680, data_out=>output_MAC_3_680);
	MAC_3_681: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_681, data_out=>output_MAC_3_681);
	MAC_3_682: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_682, data_out=>output_MAC_3_682);
	MAC_3_683: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_683, data_out=>output_MAC_3_683);
	MAC_3_684: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_684, data_out=>output_MAC_3_684);
	MAC_3_685: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_685, data_out=>output_MAC_3_685);
	MAC_3_686: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_686, data_out=>output_MAC_3_686);
	MAC_3_687: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_687, data_out=>output_MAC_3_687);
	MAC_3_688: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_688, data_out=>output_MAC_3_688);
	MAC_3_689: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_689, data_out=>output_MAC_3_689);
	MAC_3_690: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_690, data_out=>output_MAC_3_690);
	MAC_3_691: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_691, data_out=>output_MAC_3_691);
	MAC_3_692: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_692, data_out=>output_MAC_3_692);
	MAC_3_693: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_693, data_out=>output_MAC_3_693);
	MAC_3_694: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_694, data_out=>output_MAC_3_694);
	MAC_3_695: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_695, data_out=>output_MAC_3_695);
	MAC_3_696: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_696, data_out=>output_MAC_3_696);
	MAC_3_697: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_697, data_out=>output_MAC_3_697);
	MAC_3_698: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_698, data_out=>output_MAC_3_698);
	MAC_3_699: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_699, data_out=>output_MAC_3_699);
	MAC_3_700: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_700, data_out=>output_MAC_3_700);
	MAC_3_701: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_701, data_out=>output_MAC_3_701);
	MAC_3_702: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_702, data_out=>output_MAC_3_702);
	MAC_3_703: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_703, data_out=>output_MAC_3_703);
	MAC_3_704: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_704, data_out=>output_MAC_3_704);
	MAC_3_705: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_705, data_out=>output_MAC_3_705);
	MAC_3_706: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_706, data_out=>output_MAC_3_706);
	MAC_3_707: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_707, data_out=>output_MAC_3_707);
	MAC_3_708: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_708, data_out=>output_MAC_3_708);
	MAC_3_709: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_709, data_out=>output_MAC_3_709);
	MAC_3_710: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_710, data_out=>output_MAC_3_710);
	MAC_3_711: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_711, data_out=>output_MAC_3_711);
	MAC_3_712: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_712, data_out=>output_MAC_3_712);
	MAC_3_713: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_713, data_out=>output_MAC_3_713);
	MAC_3_714: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_714, data_out=>output_MAC_3_714);
	MAC_3_715: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_715, data_out=>output_MAC_3_715);
	MAC_3_716: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_716, data_out=>output_MAC_3_716);
	MAC_3_717: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_717, data_out=>output_MAC_3_717);
	MAC_3_718: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_718, data_out=>output_MAC_3_718);
	MAC_3_719: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_719, data_out=>output_MAC_3_719);
	MAC_3_720: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_720, data_out=>output_MAC_3_720);
	MAC_3_721: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_721, data_out=>output_MAC_3_721);
	MAC_3_722: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_722, data_out=>output_MAC_3_722);
	MAC_3_723: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_723, data_out=>output_MAC_3_723);
	MAC_3_724: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_724, data_out=>output_MAC_3_724);
	MAC_3_725: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_725, data_out=>output_MAC_3_725);
	MAC_3_726: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_726, data_out=>output_MAC_3_726);
	MAC_3_727: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_727, data_out=>output_MAC_3_727);
	MAC_3_728: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_728, data_out=>output_MAC_3_728);
	MAC_3_729: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_729, data_out=>output_MAC_3_729);
	MAC_3_730: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_730, data_out=>output_MAC_3_730);
	MAC_3_731: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_731, data_out=>output_MAC_3_731);
	MAC_3_732: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_732, data_out=>output_MAC_3_732);
	MAC_3_733: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_733, data_out=>output_MAC_3_733);
	MAC_3_734: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_734, data_out=>output_MAC_3_734);
	MAC_3_735: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_735, data_out=>output_MAC_3_735);
	MAC_3_736: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_736, data_out=>output_MAC_3_736);
	MAC_3_737: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_737, data_out=>output_MAC_3_737);
	MAC_3_738: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_738, data_out=>output_MAC_3_738);
	MAC_3_739: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_739, data_out=>output_MAC_3_739);
	MAC_3_740: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_740, data_out=>output_MAC_3_740);
	MAC_3_741: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_741, data_out=>output_MAC_3_741);
	MAC_3_742: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_742, data_out=>output_MAC_3_742);
	MAC_3_743: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_743, data_out=>output_MAC_3_743);
	MAC_3_744: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_744, data_out=>output_MAC_3_744);
	MAC_3_745: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_745, data_out=>output_MAC_3_745);
	MAC_3_746: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_746, data_out=>output_MAC_3_746);
	MAC_3_747: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_747, data_out=>output_MAC_3_747);
	MAC_3_748: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_748, data_out=>output_MAC_3_748);
	MAC_3_749: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_749, data_out=>output_MAC_3_749);
	MAC_3_750: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_750, data_out=>output_MAC_3_750);
	MAC_3_751: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_751, data_out=>output_MAC_3_751);
	MAC_3_752: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_752, data_out=>output_MAC_3_752);
	MAC_3_753: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_753, data_out=>output_MAC_3_753);
	MAC_3_754: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_754, data_out=>output_MAC_3_754);
	MAC_3_755: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_755, data_out=>output_MAC_3_755);
	MAC_3_756: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_756, data_out=>output_MAC_3_756);
	MAC_3_757: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_757, data_out=>output_MAC_3_757);
	MAC_3_758: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_758, data_out=>output_MAC_3_758);
	MAC_3_759: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_759, data_out=>output_MAC_3_759);
	MAC_3_760: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_760, data_out=>output_MAC_3_760);
	MAC_3_761: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_761, data_out=>output_MAC_3_761);
	MAC_3_762: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_762, data_out=>output_MAC_3_762);
	MAC_3_763: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_763, data_out=>output_MAC_3_763);
	MAC_3_764: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_764, data_out=>output_MAC_3_764);
	MAC_3_765: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_765, data_out=>output_MAC_3_765);
	MAC_3_766: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_766, data_out=>output_MAC_3_766);
	MAC_3_767: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_3, data_in_B=>input_col_767, data_out=>output_MAC_3_767);
	MAC_4_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_0, data_out=>output_MAC_4_0);
	MAC_4_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_1, data_out=>output_MAC_4_1);
	MAC_4_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_2, data_out=>output_MAC_4_2);
	MAC_4_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_3, data_out=>output_MAC_4_3);
	MAC_4_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_4, data_out=>output_MAC_4_4);
	MAC_4_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_5, data_out=>output_MAC_4_5);
	MAC_4_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_6, data_out=>output_MAC_4_6);
	MAC_4_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_7, data_out=>output_MAC_4_7);
	MAC_4_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_8, data_out=>output_MAC_4_8);
	MAC_4_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_9, data_out=>output_MAC_4_9);
	MAC_4_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_10, data_out=>output_MAC_4_10);
	MAC_4_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_11, data_out=>output_MAC_4_11);
	MAC_4_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_12, data_out=>output_MAC_4_12);
	MAC_4_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_13, data_out=>output_MAC_4_13);
	MAC_4_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_14, data_out=>output_MAC_4_14);
	MAC_4_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_15, data_out=>output_MAC_4_15);
	MAC_4_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_16, data_out=>output_MAC_4_16);
	MAC_4_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_17, data_out=>output_MAC_4_17);
	MAC_4_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_18, data_out=>output_MAC_4_18);
	MAC_4_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_19, data_out=>output_MAC_4_19);
	MAC_4_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_20, data_out=>output_MAC_4_20);
	MAC_4_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_21, data_out=>output_MAC_4_21);
	MAC_4_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_22, data_out=>output_MAC_4_22);
	MAC_4_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_23, data_out=>output_MAC_4_23);
	MAC_4_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_24, data_out=>output_MAC_4_24);
	MAC_4_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_25, data_out=>output_MAC_4_25);
	MAC_4_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_26, data_out=>output_MAC_4_26);
	MAC_4_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_27, data_out=>output_MAC_4_27);
	MAC_4_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_28, data_out=>output_MAC_4_28);
	MAC_4_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_29, data_out=>output_MAC_4_29);
	MAC_4_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_30, data_out=>output_MAC_4_30);
	MAC_4_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_31, data_out=>output_MAC_4_31);
	MAC_4_32: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_32, data_out=>output_MAC_4_32);
	MAC_4_33: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_33, data_out=>output_MAC_4_33);
	MAC_4_34: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_34, data_out=>output_MAC_4_34);
	MAC_4_35: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_35, data_out=>output_MAC_4_35);
	MAC_4_36: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_36, data_out=>output_MAC_4_36);
	MAC_4_37: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_37, data_out=>output_MAC_4_37);
	MAC_4_38: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_38, data_out=>output_MAC_4_38);
	MAC_4_39: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_39, data_out=>output_MAC_4_39);
	MAC_4_40: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_40, data_out=>output_MAC_4_40);
	MAC_4_41: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_41, data_out=>output_MAC_4_41);
	MAC_4_42: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_42, data_out=>output_MAC_4_42);
	MAC_4_43: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_43, data_out=>output_MAC_4_43);
	MAC_4_44: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_44, data_out=>output_MAC_4_44);
	MAC_4_45: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_45, data_out=>output_MAC_4_45);
	MAC_4_46: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_46, data_out=>output_MAC_4_46);
	MAC_4_47: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_47, data_out=>output_MAC_4_47);
	MAC_4_48: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_48, data_out=>output_MAC_4_48);
	MAC_4_49: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_49, data_out=>output_MAC_4_49);
	MAC_4_50: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_50, data_out=>output_MAC_4_50);
	MAC_4_51: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_51, data_out=>output_MAC_4_51);
	MAC_4_52: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_52, data_out=>output_MAC_4_52);
	MAC_4_53: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_53, data_out=>output_MAC_4_53);
	MAC_4_54: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_54, data_out=>output_MAC_4_54);
	MAC_4_55: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_55, data_out=>output_MAC_4_55);
	MAC_4_56: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_56, data_out=>output_MAC_4_56);
	MAC_4_57: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_57, data_out=>output_MAC_4_57);
	MAC_4_58: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_58, data_out=>output_MAC_4_58);
	MAC_4_59: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_59, data_out=>output_MAC_4_59);
	MAC_4_60: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_60, data_out=>output_MAC_4_60);
	MAC_4_61: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_61, data_out=>output_MAC_4_61);
	MAC_4_62: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_62, data_out=>output_MAC_4_62);
	MAC_4_63: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_63, data_out=>output_MAC_4_63);
	MAC_4_64: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_64, data_out=>output_MAC_4_64);
	MAC_4_65: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_65, data_out=>output_MAC_4_65);
	MAC_4_66: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_66, data_out=>output_MAC_4_66);
	MAC_4_67: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_67, data_out=>output_MAC_4_67);
	MAC_4_68: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_68, data_out=>output_MAC_4_68);
	MAC_4_69: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_69, data_out=>output_MAC_4_69);
	MAC_4_70: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_70, data_out=>output_MAC_4_70);
	MAC_4_71: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_71, data_out=>output_MAC_4_71);
	MAC_4_72: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_72, data_out=>output_MAC_4_72);
	MAC_4_73: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_73, data_out=>output_MAC_4_73);
	MAC_4_74: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_74, data_out=>output_MAC_4_74);
	MAC_4_75: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_75, data_out=>output_MAC_4_75);
	MAC_4_76: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_76, data_out=>output_MAC_4_76);
	MAC_4_77: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_77, data_out=>output_MAC_4_77);
	MAC_4_78: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_78, data_out=>output_MAC_4_78);
	MAC_4_79: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_79, data_out=>output_MAC_4_79);
	MAC_4_80: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_80, data_out=>output_MAC_4_80);
	MAC_4_81: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_81, data_out=>output_MAC_4_81);
	MAC_4_82: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_82, data_out=>output_MAC_4_82);
	MAC_4_83: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_83, data_out=>output_MAC_4_83);
	MAC_4_84: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_84, data_out=>output_MAC_4_84);
	MAC_4_85: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_85, data_out=>output_MAC_4_85);
	MAC_4_86: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_86, data_out=>output_MAC_4_86);
	MAC_4_87: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_87, data_out=>output_MAC_4_87);
	MAC_4_88: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_88, data_out=>output_MAC_4_88);
	MAC_4_89: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_89, data_out=>output_MAC_4_89);
	MAC_4_90: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_90, data_out=>output_MAC_4_90);
	MAC_4_91: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_91, data_out=>output_MAC_4_91);
	MAC_4_92: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_92, data_out=>output_MAC_4_92);
	MAC_4_93: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_93, data_out=>output_MAC_4_93);
	MAC_4_94: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_94, data_out=>output_MAC_4_94);
	MAC_4_95: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_95, data_out=>output_MAC_4_95);
	MAC_4_96: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_96, data_out=>output_MAC_4_96);
	MAC_4_97: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_97, data_out=>output_MAC_4_97);
	MAC_4_98: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_98, data_out=>output_MAC_4_98);
	MAC_4_99: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_99, data_out=>output_MAC_4_99);
	MAC_4_100: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_100, data_out=>output_MAC_4_100);
	MAC_4_101: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_101, data_out=>output_MAC_4_101);
	MAC_4_102: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_102, data_out=>output_MAC_4_102);
	MAC_4_103: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_103, data_out=>output_MAC_4_103);
	MAC_4_104: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_104, data_out=>output_MAC_4_104);
	MAC_4_105: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_105, data_out=>output_MAC_4_105);
	MAC_4_106: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_106, data_out=>output_MAC_4_106);
	MAC_4_107: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_107, data_out=>output_MAC_4_107);
	MAC_4_108: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_108, data_out=>output_MAC_4_108);
	MAC_4_109: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_109, data_out=>output_MAC_4_109);
	MAC_4_110: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_110, data_out=>output_MAC_4_110);
	MAC_4_111: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_111, data_out=>output_MAC_4_111);
	MAC_4_112: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_112, data_out=>output_MAC_4_112);
	MAC_4_113: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_113, data_out=>output_MAC_4_113);
	MAC_4_114: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_114, data_out=>output_MAC_4_114);
	MAC_4_115: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_115, data_out=>output_MAC_4_115);
	MAC_4_116: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_116, data_out=>output_MAC_4_116);
	MAC_4_117: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_117, data_out=>output_MAC_4_117);
	MAC_4_118: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_118, data_out=>output_MAC_4_118);
	MAC_4_119: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_119, data_out=>output_MAC_4_119);
	MAC_4_120: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_120, data_out=>output_MAC_4_120);
	MAC_4_121: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_121, data_out=>output_MAC_4_121);
	MAC_4_122: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_122, data_out=>output_MAC_4_122);
	MAC_4_123: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_123, data_out=>output_MAC_4_123);
	MAC_4_124: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_124, data_out=>output_MAC_4_124);
	MAC_4_125: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_125, data_out=>output_MAC_4_125);
	MAC_4_126: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_126, data_out=>output_MAC_4_126);
	MAC_4_127: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_127, data_out=>output_MAC_4_127);
	MAC_4_128: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_128, data_out=>output_MAC_4_128);
	MAC_4_129: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_129, data_out=>output_MAC_4_129);
	MAC_4_130: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_130, data_out=>output_MAC_4_130);
	MAC_4_131: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_131, data_out=>output_MAC_4_131);
	MAC_4_132: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_132, data_out=>output_MAC_4_132);
	MAC_4_133: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_133, data_out=>output_MAC_4_133);
	MAC_4_134: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_134, data_out=>output_MAC_4_134);
	MAC_4_135: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_135, data_out=>output_MAC_4_135);
	MAC_4_136: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_136, data_out=>output_MAC_4_136);
	MAC_4_137: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_137, data_out=>output_MAC_4_137);
	MAC_4_138: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_138, data_out=>output_MAC_4_138);
	MAC_4_139: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_139, data_out=>output_MAC_4_139);
	MAC_4_140: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_140, data_out=>output_MAC_4_140);
	MAC_4_141: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_141, data_out=>output_MAC_4_141);
	MAC_4_142: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_142, data_out=>output_MAC_4_142);
	MAC_4_143: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_143, data_out=>output_MAC_4_143);
	MAC_4_144: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_144, data_out=>output_MAC_4_144);
	MAC_4_145: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_145, data_out=>output_MAC_4_145);
	MAC_4_146: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_146, data_out=>output_MAC_4_146);
	MAC_4_147: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_147, data_out=>output_MAC_4_147);
	MAC_4_148: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_148, data_out=>output_MAC_4_148);
	MAC_4_149: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_149, data_out=>output_MAC_4_149);
	MAC_4_150: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_150, data_out=>output_MAC_4_150);
	MAC_4_151: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_151, data_out=>output_MAC_4_151);
	MAC_4_152: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_152, data_out=>output_MAC_4_152);
	MAC_4_153: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_153, data_out=>output_MAC_4_153);
	MAC_4_154: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_154, data_out=>output_MAC_4_154);
	MAC_4_155: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_155, data_out=>output_MAC_4_155);
	MAC_4_156: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_156, data_out=>output_MAC_4_156);
	MAC_4_157: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_157, data_out=>output_MAC_4_157);
	MAC_4_158: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_158, data_out=>output_MAC_4_158);
	MAC_4_159: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_159, data_out=>output_MAC_4_159);
	MAC_4_160: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_160, data_out=>output_MAC_4_160);
	MAC_4_161: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_161, data_out=>output_MAC_4_161);
	MAC_4_162: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_162, data_out=>output_MAC_4_162);
	MAC_4_163: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_163, data_out=>output_MAC_4_163);
	MAC_4_164: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_164, data_out=>output_MAC_4_164);
	MAC_4_165: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_165, data_out=>output_MAC_4_165);
	MAC_4_166: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_166, data_out=>output_MAC_4_166);
	MAC_4_167: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_167, data_out=>output_MAC_4_167);
	MAC_4_168: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_168, data_out=>output_MAC_4_168);
	MAC_4_169: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_169, data_out=>output_MAC_4_169);
	MAC_4_170: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_170, data_out=>output_MAC_4_170);
	MAC_4_171: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_171, data_out=>output_MAC_4_171);
	MAC_4_172: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_172, data_out=>output_MAC_4_172);
	MAC_4_173: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_173, data_out=>output_MAC_4_173);
	MAC_4_174: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_174, data_out=>output_MAC_4_174);
	MAC_4_175: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_175, data_out=>output_MAC_4_175);
	MAC_4_176: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_176, data_out=>output_MAC_4_176);
	MAC_4_177: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_177, data_out=>output_MAC_4_177);
	MAC_4_178: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_178, data_out=>output_MAC_4_178);
	MAC_4_179: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_179, data_out=>output_MAC_4_179);
	MAC_4_180: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_180, data_out=>output_MAC_4_180);
	MAC_4_181: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_181, data_out=>output_MAC_4_181);
	MAC_4_182: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_182, data_out=>output_MAC_4_182);
	MAC_4_183: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_183, data_out=>output_MAC_4_183);
	MAC_4_184: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_184, data_out=>output_MAC_4_184);
	MAC_4_185: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_185, data_out=>output_MAC_4_185);
	MAC_4_186: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_186, data_out=>output_MAC_4_186);
	MAC_4_187: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_187, data_out=>output_MAC_4_187);
	MAC_4_188: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_188, data_out=>output_MAC_4_188);
	MAC_4_189: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_189, data_out=>output_MAC_4_189);
	MAC_4_190: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_190, data_out=>output_MAC_4_190);
	MAC_4_191: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_191, data_out=>output_MAC_4_191);
	MAC_4_192: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_192, data_out=>output_MAC_4_192);
	MAC_4_193: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_193, data_out=>output_MAC_4_193);
	MAC_4_194: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_194, data_out=>output_MAC_4_194);
	MAC_4_195: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_195, data_out=>output_MAC_4_195);
	MAC_4_196: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_196, data_out=>output_MAC_4_196);
	MAC_4_197: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_197, data_out=>output_MAC_4_197);
	MAC_4_198: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_198, data_out=>output_MAC_4_198);
	MAC_4_199: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_199, data_out=>output_MAC_4_199);
	MAC_4_200: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_200, data_out=>output_MAC_4_200);
	MAC_4_201: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_201, data_out=>output_MAC_4_201);
	MAC_4_202: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_202, data_out=>output_MAC_4_202);
	MAC_4_203: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_203, data_out=>output_MAC_4_203);
	MAC_4_204: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_204, data_out=>output_MAC_4_204);
	MAC_4_205: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_205, data_out=>output_MAC_4_205);
	MAC_4_206: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_206, data_out=>output_MAC_4_206);
	MAC_4_207: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_207, data_out=>output_MAC_4_207);
	MAC_4_208: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_208, data_out=>output_MAC_4_208);
	MAC_4_209: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_209, data_out=>output_MAC_4_209);
	MAC_4_210: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_210, data_out=>output_MAC_4_210);
	MAC_4_211: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_211, data_out=>output_MAC_4_211);
	MAC_4_212: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_212, data_out=>output_MAC_4_212);
	MAC_4_213: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_213, data_out=>output_MAC_4_213);
	MAC_4_214: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_214, data_out=>output_MAC_4_214);
	MAC_4_215: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_215, data_out=>output_MAC_4_215);
	MAC_4_216: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_216, data_out=>output_MAC_4_216);
	MAC_4_217: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_217, data_out=>output_MAC_4_217);
	MAC_4_218: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_218, data_out=>output_MAC_4_218);
	MAC_4_219: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_219, data_out=>output_MAC_4_219);
	MAC_4_220: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_220, data_out=>output_MAC_4_220);
	MAC_4_221: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_221, data_out=>output_MAC_4_221);
	MAC_4_222: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_222, data_out=>output_MAC_4_222);
	MAC_4_223: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_223, data_out=>output_MAC_4_223);
	MAC_4_224: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_224, data_out=>output_MAC_4_224);
	MAC_4_225: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_225, data_out=>output_MAC_4_225);
	MAC_4_226: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_226, data_out=>output_MAC_4_226);
	MAC_4_227: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_227, data_out=>output_MAC_4_227);
	MAC_4_228: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_228, data_out=>output_MAC_4_228);
	MAC_4_229: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_229, data_out=>output_MAC_4_229);
	MAC_4_230: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_230, data_out=>output_MAC_4_230);
	MAC_4_231: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_231, data_out=>output_MAC_4_231);
	MAC_4_232: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_232, data_out=>output_MAC_4_232);
	MAC_4_233: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_233, data_out=>output_MAC_4_233);
	MAC_4_234: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_234, data_out=>output_MAC_4_234);
	MAC_4_235: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_235, data_out=>output_MAC_4_235);
	MAC_4_236: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_236, data_out=>output_MAC_4_236);
	MAC_4_237: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_237, data_out=>output_MAC_4_237);
	MAC_4_238: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_238, data_out=>output_MAC_4_238);
	MAC_4_239: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_239, data_out=>output_MAC_4_239);
	MAC_4_240: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_240, data_out=>output_MAC_4_240);
	MAC_4_241: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_241, data_out=>output_MAC_4_241);
	MAC_4_242: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_242, data_out=>output_MAC_4_242);
	MAC_4_243: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_243, data_out=>output_MAC_4_243);
	MAC_4_244: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_244, data_out=>output_MAC_4_244);
	MAC_4_245: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_245, data_out=>output_MAC_4_245);
	MAC_4_246: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_246, data_out=>output_MAC_4_246);
	MAC_4_247: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_247, data_out=>output_MAC_4_247);
	MAC_4_248: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_248, data_out=>output_MAC_4_248);
	MAC_4_249: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_249, data_out=>output_MAC_4_249);
	MAC_4_250: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_250, data_out=>output_MAC_4_250);
	MAC_4_251: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_251, data_out=>output_MAC_4_251);
	MAC_4_252: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_252, data_out=>output_MAC_4_252);
	MAC_4_253: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_253, data_out=>output_MAC_4_253);
	MAC_4_254: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_254, data_out=>output_MAC_4_254);
	MAC_4_255: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_255, data_out=>output_MAC_4_255);
	MAC_4_256: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_256, data_out=>output_MAC_4_256);
	MAC_4_257: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_257, data_out=>output_MAC_4_257);
	MAC_4_258: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_258, data_out=>output_MAC_4_258);
	MAC_4_259: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_259, data_out=>output_MAC_4_259);
	MAC_4_260: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_260, data_out=>output_MAC_4_260);
	MAC_4_261: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_261, data_out=>output_MAC_4_261);
	MAC_4_262: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_262, data_out=>output_MAC_4_262);
	MAC_4_263: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_263, data_out=>output_MAC_4_263);
	MAC_4_264: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_264, data_out=>output_MAC_4_264);
	MAC_4_265: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_265, data_out=>output_MAC_4_265);
	MAC_4_266: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_266, data_out=>output_MAC_4_266);
	MAC_4_267: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_267, data_out=>output_MAC_4_267);
	MAC_4_268: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_268, data_out=>output_MAC_4_268);
	MAC_4_269: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_269, data_out=>output_MAC_4_269);
	MAC_4_270: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_270, data_out=>output_MAC_4_270);
	MAC_4_271: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_271, data_out=>output_MAC_4_271);
	MAC_4_272: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_272, data_out=>output_MAC_4_272);
	MAC_4_273: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_273, data_out=>output_MAC_4_273);
	MAC_4_274: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_274, data_out=>output_MAC_4_274);
	MAC_4_275: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_275, data_out=>output_MAC_4_275);
	MAC_4_276: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_276, data_out=>output_MAC_4_276);
	MAC_4_277: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_277, data_out=>output_MAC_4_277);
	MAC_4_278: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_278, data_out=>output_MAC_4_278);
	MAC_4_279: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_279, data_out=>output_MAC_4_279);
	MAC_4_280: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_280, data_out=>output_MAC_4_280);
	MAC_4_281: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_281, data_out=>output_MAC_4_281);
	MAC_4_282: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_282, data_out=>output_MAC_4_282);
	MAC_4_283: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_283, data_out=>output_MAC_4_283);
	MAC_4_284: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_284, data_out=>output_MAC_4_284);
	MAC_4_285: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_285, data_out=>output_MAC_4_285);
	MAC_4_286: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_286, data_out=>output_MAC_4_286);
	MAC_4_287: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_287, data_out=>output_MAC_4_287);
	MAC_4_288: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_288, data_out=>output_MAC_4_288);
	MAC_4_289: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_289, data_out=>output_MAC_4_289);
	MAC_4_290: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_290, data_out=>output_MAC_4_290);
	MAC_4_291: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_291, data_out=>output_MAC_4_291);
	MAC_4_292: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_292, data_out=>output_MAC_4_292);
	MAC_4_293: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_293, data_out=>output_MAC_4_293);
	MAC_4_294: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_294, data_out=>output_MAC_4_294);
	MAC_4_295: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_295, data_out=>output_MAC_4_295);
	MAC_4_296: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_296, data_out=>output_MAC_4_296);
	MAC_4_297: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_297, data_out=>output_MAC_4_297);
	MAC_4_298: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_298, data_out=>output_MAC_4_298);
	MAC_4_299: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_299, data_out=>output_MAC_4_299);
	MAC_4_300: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_300, data_out=>output_MAC_4_300);
	MAC_4_301: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_301, data_out=>output_MAC_4_301);
	MAC_4_302: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_302, data_out=>output_MAC_4_302);
	MAC_4_303: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_303, data_out=>output_MAC_4_303);
	MAC_4_304: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_304, data_out=>output_MAC_4_304);
	MAC_4_305: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_305, data_out=>output_MAC_4_305);
	MAC_4_306: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_306, data_out=>output_MAC_4_306);
	MAC_4_307: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_307, data_out=>output_MAC_4_307);
	MAC_4_308: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_308, data_out=>output_MAC_4_308);
	MAC_4_309: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_309, data_out=>output_MAC_4_309);
	MAC_4_310: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_310, data_out=>output_MAC_4_310);
	MAC_4_311: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_311, data_out=>output_MAC_4_311);
	MAC_4_312: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_312, data_out=>output_MAC_4_312);
	MAC_4_313: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_313, data_out=>output_MAC_4_313);
	MAC_4_314: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_314, data_out=>output_MAC_4_314);
	MAC_4_315: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_315, data_out=>output_MAC_4_315);
	MAC_4_316: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_316, data_out=>output_MAC_4_316);
	MAC_4_317: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_317, data_out=>output_MAC_4_317);
	MAC_4_318: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_318, data_out=>output_MAC_4_318);
	MAC_4_319: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_319, data_out=>output_MAC_4_319);
	MAC_4_320: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_320, data_out=>output_MAC_4_320);
	MAC_4_321: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_321, data_out=>output_MAC_4_321);
	MAC_4_322: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_322, data_out=>output_MAC_4_322);
	MAC_4_323: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_323, data_out=>output_MAC_4_323);
	MAC_4_324: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_324, data_out=>output_MAC_4_324);
	MAC_4_325: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_325, data_out=>output_MAC_4_325);
	MAC_4_326: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_326, data_out=>output_MAC_4_326);
	MAC_4_327: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_327, data_out=>output_MAC_4_327);
	MAC_4_328: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_328, data_out=>output_MAC_4_328);
	MAC_4_329: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_329, data_out=>output_MAC_4_329);
	MAC_4_330: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_330, data_out=>output_MAC_4_330);
	MAC_4_331: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_331, data_out=>output_MAC_4_331);
	MAC_4_332: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_332, data_out=>output_MAC_4_332);
	MAC_4_333: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_333, data_out=>output_MAC_4_333);
	MAC_4_334: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_334, data_out=>output_MAC_4_334);
	MAC_4_335: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_335, data_out=>output_MAC_4_335);
	MAC_4_336: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_336, data_out=>output_MAC_4_336);
	MAC_4_337: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_337, data_out=>output_MAC_4_337);
	MAC_4_338: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_338, data_out=>output_MAC_4_338);
	MAC_4_339: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_339, data_out=>output_MAC_4_339);
	MAC_4_340: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_340, data_out=>output_MAC_4_340);
	MAC_4_341: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_341, data_out=>output_MAC_4_341);
	MAC_4_342: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_342, data_out=>output_MAC_4_342);
	MAC_4_343: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_343, data_out=>output_MAC_4_343);
	MAC_4_344: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_344, data_out=>output_MAC_4_344);
	MAC_4_345: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_345, data_out=>output_MAC_4_345);
	MAC_4_346: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_346, data_out=>output_MAC_4_346);
	MAC_4_347: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_347, data_out=>output_MAC_4_347);
	MAC_4_348: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_348, data_out=>output_MAC_4_348);
	MAC_4_349: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_349, data_out=>output_MAC_4_349);
	MAC_4_350: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_350, data_out=>output_MAC_4_350);
	MAC_4_351: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_351, data_out=>output_MAC_4_351);
	MAC_4_352: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_352, data_out=>output_MAC_4_352);
	MAC_4_353: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_353, data_out=>output_MAC_4_353);
	MAC_4_354: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_354, data_out=>output_MAC_4_354);
	MAC_4_355: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_355, data_out=>output_MAC_4_355);
	MAC_4_356: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_356, data_out=>output_MAC_4_356);
	MAC_4_357: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_357, data_out=>output_MAC_4_357);
	MAC_4_358: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_358, data_out=>output_MAC_4_358);
	MAC_4_359: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_359, data_out=>output_MAC_4_359);
	MAC_4_360: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_360, data_out=>output_MAC_4_360);
	MAC_4_361: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_361, data_out=>output_MAC_4_361);
	MAC_4_362: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_362, data_out=>output_MAC_4_362);
	MAC_4_363: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_363, data_out=>output_MAC_4_363);
	MAC_4_364: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_364, data_out=>output_MAC_4_364);
	MAC_4_365: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_365, data_out=>output_MAC_4_365);
	MAC_4_366: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_366, data_out=>output_MAC_4_366);
	MAC_4_367: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_367, data_out=>output_MAC_4_367);
	MAC_4_368: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_368, data_out=>output_MAC_4_368);
	MAC_4_369: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_369, data_out=>output_MAC_4_369);
	MAC_4_370: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_370, data_out=>output_MAC_4_370);
	MAC_4_371: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_371, data_out=>output_MAC_4_371);
	MAC_4_372: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_372, data_out=>output_MAC_4_372);
	MAC_4_373: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_373, data_out=>output_MAC_4_373);
	MAC_4_374: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_374, data_out=>output_MAC_4_374);
	MAC_4_375: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_375, data_out=>output_MAC_4_375);
	MAC_4_376: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_376, data_out=>output_MAC_4_376);
	MAC_4_377: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_377, data_out=>output_MAC_4_377);
	MAC_4_378: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_378, data_out=>output_MAC_4_378);
	MAC_4_379: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_379, data_out=>output_MAC_4_379);
	MAC_4_380: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_380, data_out=>output_MAC_4_380);
	MAC_4_381: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_381, data_out=>output_MAC_4_381);
	MAC_4_382: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_382, data_out=>output_MAC_4_382);
	MAC_4_383: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_383, data_out=>output_MAC_4_383);
	MAC_4_384: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_384, data_out=>output_MAC_4_384);
	MAC_4_385: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_385, data_out=>output_MAC_4_385);
	MAC_4_386: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_386, data_out=>output_MAC_4_386);
	MAC_4_387: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_387, data_out=>output_MAC_4_387);
	MAC_4_388: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_388, data_out=>output_MAC_4_388);
	MAC_4_389: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_389, data_out=>output_MAC_4_389);
	MAC_4_390: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_390, data_out=>output_MAC_4_390);
	MAC_4_391: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_391, data_out=>output_MAC_4_391);
	MAC_4_392: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_392, data_out=>output_MAC_4_392);
	MAC_4_393: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_393, data_out=>output_MAC_4_393);
	MAC_4_394: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_394, data_out=>output_MAC_4_394);
	MAC_4_395: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_395, data_out=>output_MAC_4_395);
	MAC_4_396: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_396, data_out=>output_MAC_4_396);
	MAC_4_397: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_397, data_out=>output_MAC_4_397);
	MAC_4_398: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_398, data_out=>output_MAC_4_398);
	MAC_4_399: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_399, data_out=>output_MAC_4_399);
	MAC_4_400: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_400, data_out=>output_MAC_4_400);
	MAC_4_401: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_401, data_out=>output_MAC_4_401);
	MAC_4_402: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_402, data_out=>output_MAC_4_402);
	MAC_4_403: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_403, data_out=>output_MAC_4_403);
	MAC_4_404: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_404, data_out=>output_MAC_4_404);
	MAC_4_405: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_405, data_out=>output_MAC_4_405);
	MAC_4_406: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_406, data_out=>output_MAC_4_406);
	MAC_4_407: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_407, data_out=>output_MAC_4_407);
	MAC_4_408: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_408, data_out=>output_MAC_4_408);
	MAC_4_409: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_409, data_out=>output_MAC_4_409);
	MAC_4_410: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_410, data_out=>output_MAC_4_410);
	MAC_4_411: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_411, data_out=>output_MAC_4_411);
	MAC_4_412: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_412, data_out=>output_MAC_4_412);
	MAC_4_413: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_413, data_out=>output_MAC_4_413);
	MAC_4_414: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_414, data_out=>output_MAC_4_414);
	MAC_4_415: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_415, data_out=>output_MAC_4_415);
	MAC_4_416: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_416, data_out=>output_MAC_4_416);
	MAC_4_417: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_417, data_out=>output_MAC_4_417);
	MAC_4_418: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_418, data_out=>output_MAC_4_418);
	MAC_4_419: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_419, data_out=>output_MAC_4_419);
	MAC_4_420: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_420, data_out=>output_MAC_4_420);
	MAC_4_421: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_421, data_out=>output_MAC_4_421);
	MAC_4_422: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_422, data_out=>output_MAC_4_422);
	MAC_4_423: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_423, data_out=>output_MAC_4_423);
	MAC_4_424: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_424, data_out=>output_MAC_4_424);
	MAC_4_425: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_425, data_out=>output_MAC_4_425);
	MAC_4_426: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_426, data_out=>output_MAC_4_426);
	MAC_4_427: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_427, data_out=>output_MAC_4_427);
	MAC_4_428: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_428, data_out=>output_MAC_4_428);
	MAC_4_429: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_429, data_out=>output_MAC_4_429);
	MAC_4_430: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_430, data_out=>output_MAC_4_430);
	MAC_4_431: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_431, data_out=>output_MAC_4_431);
	MAC_4_432: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_432, data_out=>output_MAC_4_432);
	MAC_4_433: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_433, data_out=>output_MAC_4_433);
	MAC_4_434: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_434, data_out=>output_MAC_4_434);
	MAC_4_435: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_435, data_out=>output_MAC_4_435);
	MAC_4_436: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_436, data_out=>output_MAC_4_436);
	MAC_4_437: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_437, data_out=>output_MAC_4_437);
	MAC_4_438: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_438, data_out=>output_MAC_4_438);
	MAC_4_439: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_439, data_out=>output_MAC_4_439);
	MAC_4_440: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_440, data_out=>output_MAC_4_440);
	MAC_4_441: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_441, data_out=>output_MAC_4_441);
	MAC_4_442: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_442, data_out=>output_MAC_4_442);
	MAC_4_443: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_443, data_out=>output_MAC_4_443);
	MAC_4_444: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_444, data_out=>output_MAC_4_444);
	MAC_4_445: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_445, data_out=>output_MAC_4_445);
	MAC_4_446: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_446, data_out=>output_MAC_4_446);
	MAC_4_447: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_447, data_out=>output_MAC_4_447);
	MAC_4_448: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_448, data_out=>output_MAC_4_448);
	MAC_4_449: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_449, data_out=>output_MAC_4_449);
	MAC_4_450: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_450, data_out=>output_MAC_4_450);
	MAC_4_451: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_451, data_out=>output_MAC_4_451);
	MAC_4_452: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_452, data_out=>output_MAC_4_452);
	MAC_4_453: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_453, data_out=>output_MAC_4_453);
	MAC_4_454: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_454, data_out=>output_MAC_4_454);
	MAC_4_455: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_455, data_out=>output_MAC_4_455);
	MAC_4_456: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_456, data_out=>output_MAC_4_456);
	MAC_4_457: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_457, data_out=>output_MAC_4_457);
	MAC_4_458: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_458, data_out=>output_MAC_4_458);
	MAC_4_459: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_459, data_out=>output_MAC_4_459);
	MAC_4_460: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_460, data_out=>output_MAC_4_460);
	MAC_4_461: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_461, data_out=>output_MAC_4_461);
	MAC_4_462: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_462, data_out=>output_MAC_4_462);
	MAC_4_463: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_463, data_out=>output_MAC_4_463);
	MAC_4_464: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_464, data_out=>output_MAC_4_464);
	MAC_4_465: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_465, data_out=>output_MAC_4_465);
	MAC_4_466: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_466, data_out=>output_MAC_4_466);
	MAC_4_467: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_467, data_out=>output_MAC_4_467);
	MAC_4_468: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_468, data_out=>output_MAC_4_468);
	MAC_4_469: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_469, data_out=>output_MAC_4_469);
	MAC_4_470: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_470, data_out=>output_MAC_4_470);
	MAC_4_471: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_471, data_out=>output_MAC_4_471);
	MAC_4_472: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_472, data_out=>output_MAC_4_472);
	MAC_4_473: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_473, data_out=>output_MAC_4_473);
	MAC_4_474: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_474, data_out=>output_MAC_4_474);
	MAC_4_475: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_475, data_out=>output_MAC_4_475);
	MAC_4_476: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_476, data_out=>output_MAC_4_476);
	MAC_4_477: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_477, data_out=>output_MAC_4_477);
	MAC_4_478: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_478, data_out=>output_MAC_4_478);
	MAC_4_479: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_479, data_out=>output_MAC_4_479);
	MAC_4_480: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_480, data_out=>output_MAC_4_480);
	MAC_4_481: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_481, data_out=>output_MAC_4_481);
	MAC_4_482: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_482, data_out=>output_MAC_4_482);
	MAC_4_483: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_483, data_out=>output_MAC_4_483);
	MAC_4_484: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_484, data_out=>output_MAC_4_484);
	MAC_4_485: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_485, data_out=>output_MAC_4_485);
	MAC_4_486: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_486, data_out=>output_MAC_4_486);
	MAC_4_487: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_487, data_out=>output_MAC_4_487);
	MAC_4_488: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_488, data_out=>output_MAC_4_488);
	MAC_4_489: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_489, data_out=>output_MAC_4_489);
	MAC_4_490: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_490, data_out=>output_MAC_4_490);
	MAC_4_491: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_491, data_out=>output_MAC_4_491);
	MAC_4_492: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_492, data_out=>output_MAC_4_492);
	MAC_4_493: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_493, data_out=>output_MAC_4_493);
	MAC_4_494: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_494, data_out=>output_MAC_4_494);
	MAC_4_495: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_495, data_out=>output_MAC_4_495);
	MAC_4_496: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_496, data_out=>output_MAC_4_496);
	MAC_4_497: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_497, data_out=>output_MAC_4_497);
	MAC_4_498: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_498, data_out=>output_MAC_4_498);
	MAC_4_499: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_499, data_out=>output_MAC_4_499);
	MAC_4_500: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_500, data_out=>output_MAC_4_500);
	MAC_4_501: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_501, data_out=>output_MAC_4_501);
	MAC_4_502: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_502, data_out=>output_MAC_4_502);
	MAC_4_503: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_503, data_out=>output_MAC_4_503);
	MAC_4_504: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_504, data_out=>output_MAC_4_504);
	MAC_4_505: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_505, data_out=>output_MAC_4_505);
	MAC_4_506: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_506, data_out=>output_MAC_4_506);
	MAC_4_507: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_507, data_out=>output_MAC_4_507);
	MAC_4_508: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_508, data_out=>output_MAC_4_508);
	MAC_4_509: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_509, data_out=>output_MAC_4_509);
	MAC_4_510: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_510, data_out=>output_MAC_4_510);
	MAC_4_511: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_511, data_out=>output_MAC_4_511);
	MAC_4_512: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_512, data_out=>output_MAC_4_512);
	MAC_4_513: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_513, data_out=>output_MAC_4_513);
	MAC_4_514: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_514, data_out=>output_MAC_4_514);
	MAC_4_515: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_515, data_out=>output_MAC_4_515);
	MAC_4_516: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_516, data_out=>output_MAC_4_516);
	MAC_4_517: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_517, data_out=>output_MAC_4_517);
	MAC_4_518: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_518, data_out=>output_MAC_4_518);
	MAC_4_519: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_519, data_out=>output_MAC_4_519);
	MAC_4_520: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_520, data_out=>output_MAC_4_520);
	MAC_4_521: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_521, data_out=>output_MAC_4_521);
	MAC_4_522: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_522, data_out=>output_MAC_4_522);
	MAC_4_523: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_523, data_out=>output_MAC_4_523);
	MAC_4_524: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_524, data_out=>output_MAC_4_524);
	MAC_4_525: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_525, data_out=>output_MAC_4_525);
	MAC_4_526: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_526, data_out=>output_MAC_4_526);
	MAC_4_527: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_527, data_out=>output_MAC_4_527);
	MAC_4_528: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_528, data_out=>output_MAC_4_528);
	MAC_4_529: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_529, data_out=>output_MAC_4_529);
	MAC_4_530: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_530, data_out=>output_MAC_4_530);
	MAC_4_531: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_531, data_out=>output_MAC_4_531);
	MAC_4_532: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_532, data_out=>output_MAC_4_532);
	MAC_4_533: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_533, data_out=>output_MAC_4_533);
	MAC_4_534: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_534, data_out=>output_MAC_4_534);
	MAC_4_535: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_535, data_out=>output_MAC_4_535);
	MAC_4_536: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_536, data_out=>output_MAC_4_536);
	MAC_4_537: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_537, data_out=>output_MAC_4_537);
	MAC_4_538: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_538, data_out=>output_MAC_4_538);
	MAC_4_539: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_539, data_out=>output_MAC_4_539);
	MAC_4_540: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_540, data_out=>output_MAC_4_540);
	MAC_4_541: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_541, data_out=>output_MAC_4_541);
	MAC_4_542: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_542, data_out=>output_MAC_4_542);
	MAC_4_543: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_543, data_out=>output_MAC_4_543);
	MAC_4_544: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_544, data_out=>output_MAC_4_544);
	MAC_4_545: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_545, data_out=>output_MAC_4_545);
	MAC_4_546: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_546, data_out=>output_MAC_4_546);
	MAC_4_547: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_547, data_out=>output_MAC_4_547);
	MAC_4_548: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_548, data_out=>output_MAC_4_548);
	MAC_4_549: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_549, data_out=>output_MAC_4_549);
	MAC_4_550: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_550, data_out=>output_MAC_4_550);
	MAC_4_551: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_551, data_out=>output_MAC_4_551);
	MAC_4_552: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_552, data_out=>output_MAC_4_552);
	MAC_4_553: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_553, data_out=>output_MAC_4_553);
	MAC_4_554: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_554, data_out=>output_MAC_4_554);
	MAC_4_555: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_555, data_out=>output_MAC_4_555);
	MAC_4_556: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_556, data_out=>output_MAC_4_556);
	MAC_4_557: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_557, data_out=>output_MAC_4_557);
	MAC_4_558: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_558, data_out=>output_MAC_4_558);
	MAC_4_559: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_559, data_out=>output_MAC_4_559);
	MAC_4_560: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_560, data_out=>output_MAC_4_560);
	MAC_4_561: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_561, data_out=>output_MAC_4_561);
	MAC_4_562: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_562, data_out=>output_MAC_4_562);
	MAC_4_563: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_563, data_out=>output_MAC_4_563);
	MAC_4_564: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_564, data_out=>output_MAC_4_564);
	MAC_4_565: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_565, data_out=>output_MAC_4_565);
	MAC_4_566: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_566, data_out=>output_MAC_4_566);
	MAC_4_567: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_567, data_out=>output_MAC_4_567);
	MAC_4_568: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_568, data_out=>output_MAC_4_568);
	MAC_4_569: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_569, data_out=>output_MAC_4_569);
	MAC_4_570: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_570, data_out=>output_MAC_4_570);
	MAC_4_571: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_571, data_out=>output_MAC_4_571);
	MAC_4_572: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_572, data_out=>output_MAC_4_572);
	MAC_4_573: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_573, data_out=>output_MAC_4_573);
	MAC_4_574: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_574, data_out=>output_MAC_4_574);
	MAC_4_575: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_575, data_out=>output_MAC_4_575);
	MAC_4_576: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_576, data_out=>output_MAC_4_576);
	MAC_4_577: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_577, data_out=>output_MAC_4_577);
	MAC_4_578: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_578, data_out=>output_MAC_4_578);
	MAC_4_579: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_579, data_out=>output_MAC_4_579);
	MAC_4_580: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_580, data_out=>output_MAC_4_580);
	MAC_4_581: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_581, data_out=>output_MAC_4_581);
	MAC_4_582: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_582, data_out=>output_MAC_4_582);
	MAC_4_583: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_583, data_out=>output_MAC_4_583);
	MAC_4_584: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_584, data_out=>output_MAC_4_584);
	MAC_4_585: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_585, data_out=>output_MAC_4_585);
	MAC_4_586: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_586, data_out=>output_MAC_4_586);
	MAC_4_587: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_587, data_out=>output_MAC_4_587);
	MAC_4_588: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_588, data_out=>output_MAC_4_588);
	MAC_4_589: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_589, data_out=>output_MAC_4_589);
	MAC_4_590: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_590, data_out=>output_MAC_4_590);
	MAC_4_591: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_591, data_out=>output_MAC_4_591);
	MAC_4_592: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_592, data_out=>output_MAC_4_592);
	MAC_4_593: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_593, data_out=>output_MAC_4_593);
	MAC_4_594: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_594, data_out=>output_MAC_4_594);
	MAC_4_595: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_595, data_out=>output_MAC_4_595);
	MAC_4_596: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_596, data_out=>output_MAC_4_596);
	MAC_4_597: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_597, data_out=>output_MAC_4_597);
	MAC_4_598: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_598, data_out=>output_MAC_4_598);
	MAC_4_599: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_599, data_out=>output_MAC_4_599);
	MAC_4_600: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_600, data_out=>output_MAC_4_600);
	MAC_4_601: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_601, data_out=>output_MAC_4_601);
	MAC_4_602: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_602, data_out=>output_MAC_4_602);
	MAC_4_603: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_603, data_out=>output_MAC_4_603);
	MAC_4_604: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_604, data_out=>output_MAC_4_604);
	MAC_4_605: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_605, data_out=>output_MAC_4_605);
	MAC_4_606: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_606, data_out=>output_MAC_4_606);
	MAC_4_607: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_607, data_out=>output_MAC_4_607);
	MAC_4_608: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_608, data_out=>output_MAC_4_608);
	MAC_4_609: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_609, data_out=>output_MAC_4_609);
	MAC_4_610: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_610, data_out=>output_MAC_4_610);
	MAC_4_611: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_611, data_out=>output_MAC_4_611);
	MAC_4_612: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_612, data_out=>output_MAC_4_612);
	MAC_4_613: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_613, data_out=>output_MAC_4_613);
	MAC_4_614: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_614, data_out=>output_MAC_4_614);
	MAC_4_615: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_615, data_out=>output_MAC_4_615);
	MAC_4_616: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_616, data_out=>output_MAC_4_616);
	MAC_4_617: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_617, data_out=>output_MAC_4_617);
	MAC_4_618: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_618, data_out=>output_MAC_4_618);
	MAC_4_619: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_619, data_out=>output_MAC_4_619);
	MAC_4_620: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_620, data_out=>output_MAC_4_620);
	MAC_4_621: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_621, data_out=>output_MAC_4_621);
	MAC_4_622: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_622, data_out=>output_MAC_4_622);
	MAC_4_623: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_623, data_out=>output_MAC_4_623);
	MAC_4_624: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_624, data_out=>output_MAC_4_624);
	MAC_4_625: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_625, data_out=>output_MAC_4_625);
	MAC_4_626: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_626, data_out=>output_MAC_4_626);
	MAC_4_627: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_627, data_out=>output_MAC_4_627);
	MAC_4_628: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_628, data_out=>output_MAC_4_628);
	MAC_4_629: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_629, data_out=>output_MAC_4_629);
	MAC_4_630: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_630, data_out=>output_MAC_4_630);
	MAC_4_631: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_631, data_out=>output_MAC_4_631);
	MAC_4_632: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_632, data_out=>output_MAC_4_632);
	MAC_4_633: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_633, data_out=>output_MAC_4_633);
	MAC_4_634: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_634, data_out=>output_MAC_4_634);
	MAC_4_635: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_635, data_out=>output_MAC_4_635);
	MAC_4_636: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_636, data_out=>output_MAC_4_636);
	MAC_4_637: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_637, data_out=>output_MAC_4_637);
	MAC_4_638: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_638, data_out=>output_MAC_4_638);
	MAC_4_639: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_639, data_out=>output_MAC_4_639);
	MAC_4_640: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_640, data_out=>output_MAC_4_640);
	MAC_4_641: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_641, data_out=>output_MAC_4_641);
	MAC_4_642: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_642, data_out=>output_MAC_4_642);
	MAC_4_643: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_643, data_out=>output_MAC_4_643);
	MAC_4_644: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_644, data_out=>output_MAC_4_644);
	MAC_4_645: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_645, data_out=>output_MAC_4_645);
	MAC_4_646: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_646, data_out=>output_MAC_4_646);
	MAC_4_647: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_647, data_out=>output_MAC_4_647);
	MAC_4_648: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_648, data_out=>output_MAC_4_648);
	MAC_4_649: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_649, data_out=>output_MAC_4_649);
	MAC_4_650: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_650, data_out=>output_MAC_4_650);
	MAC_4_651: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_651, data_out=>output_MAC_4_651);
	MAC_4_652: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_652, data_out=>output_MAC_4_652);
	MAC_4_653: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_653, data_out=>output_MAC_4_653);
	MAC_4_654: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_654, data_out=>output_MAC_4_654);
	MAC_4_655: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_655, data_out=>output_MAC_4_655);
	MAC_4_656: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_656, data_out=>output_MAC_4_656);
	MAC_4_657: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_657, data_out=>output_MAC_4_657);
	MAC_4_658: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_658, data_out=>output_MAC_4_658);
	MAC_4_659: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_659, data_out=>output_MAC_4_659);
	MAC_4_660: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_660, data_out=>output_MAC_4_660);
	MAC_4_661: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_661, data_out=>output_MAC_4_661);
	MAC_4_662: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_662, data_out=>output_MAC_4_662);
	MAC_4_663: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_663, data_out=>output_MAC_4_663);
	MAC_4_664: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_664, data_out=>output_MAC_4_664);
	MAC_4_665: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_665, data_out=>output_MAC_4_665);
	MAC_4_666: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_666, data_out=>output_MAC_4_666);
	MAC_4_667: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_667, data_out=>output_MAC_4_667);
	MAC_4_668: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_668, data_out=>output_MAC_4_668);
	MAC_4_669: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_669, data_out=>output_MAC_4_669);
	MAC_4_670: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_670, data_out=>output_MAC_4_670);
	MAC_4_671: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_671, data_out=>output_MAC_4_671);
	MAC_4_672: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_672, data_out=>output_MAC_4_672);
	MAC_4_673: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_673, data_out=>output_MAC_4_673);
	MAC_4_674: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_674, data_out=>output_MAC_4_674);
	MAC_4_675: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_675, data_out=>output_MAC_4_675);
	MAC_4_676: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_676, data_out=>output_MAC_4_676);
	MAC_4_677: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_677, data_out=>output_MAC_4_677);
	MAC_4_678: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_678, data_out=>output_MAC_4_678);
	MAC_4_679: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_679, data_out=>output_MAC_4_679);
	MAC_4_680: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_680, data_out=>output_MAC_4_680);
	MAC_4_681: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_681, data_out=>output_MAC_4_681);
	MAC_4_682: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_682, data_out=>output_MAC_4_682);
	MAC_4_683: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_683, data_out=>output_MAC_4_683);
	MAC_4_684: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_684, data_out=>output_MAC_4_684);
	MAC_4_685: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_685, data_out=>output_MAC_4_685);
	MAC_4_686: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_686, data_out=>output_MAC_4_686);
	MAC_4_687: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_687, data_out=>output_MAC_4_687);
	MAC_4_688: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_688, data_out=>output_MAC_4_688);
	MAC_4_689: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_689, data_out=>output_MAC_4_689);
	MAC_4_690: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_690, data_out=>output_MAC_4_690);
	MAC_4_691: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_691, data_out=>output_MAC_4_691);
	MAC_4_692: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_692, data_out=>output_MAC_4_692);
	MAC_4_693: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_693, data_out=>output_MAC_4_693);
	MAC_4_694: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_694, data_out=>output_MAC_4_694);
	MAC_4_695: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_695, data_out=>output_MAC_4_695);
	MAC_4_696: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_696, data_out=>output_MAC_4_696);
	MAC_4_697: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_697, data_out=>output_MAC_4_697);
	MAC_4_698: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_698, data_out=>output_MAC_4_698);
	MAC_4_699: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_699, data_out=>output_MAC_4_699);
	MAC_4_700: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_700, data_out=>output_MAC_4_700);
	MAC_4_701: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_701, data_out=>output_MAC_4_701);
	MAC_4_702: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_702, data_out=>output_MAC_4_702);
	MAC_4_703: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_703, data_out=>output_MAC_4_703);
	MAC_4_704: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_704, data_out=>output_MAC_4_704);
	MAC_4_705: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_705, data_out=>output_MAC_4_705);
	MAC_4_706: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_706, data_out=>output_MAC_4_706);
	MAC_4_707: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_707, data_out=>output_MAC_4_707);
	MAC_4_708: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_708, data_out=>output_MAC_4_708);
	MAC_4_709: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_709, data_out=>output_MAC_4_709);
	MAC_4_710: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_710, data_out=>output_MAC_4_710);
	MAC_4_711: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_711, data_out=>output_MAC_4_711);
	MAC_4_712: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_712, data_out=>output_MAC_4_712);
	MAC_4_713: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_713, data_out=>output_MAC_4_713);
	MAC_4_714: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_714, data_out=>output_MAC_4_714);
	MAC_4_715: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_715, data_out=>output_MAC_4_715);
	MAC_4_716: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_716, data_out=>output_MAC_4_716);
	MAC_4_717: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_717, data_out=>output_MAC_4_717);
	MAC_4_718: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_718, data_out=>output_MAC_4_718);
	MAC_4_719: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_719, data_out=>output_MAC_4_719);
	MAC_4_720: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_720, data_out=>output_MAC_4_720);
	MAC_4_721: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_721, data_out=>output_MAC_4_721);
	MAC_4_722: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_722, data_out=>output_MAC_4_722);
	MAC_4_723: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_723, data_out=>output_MAC_4_723);
	MAC_4_724: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_724, data_out=>output_MAC_4_724);
	MAC_4_725: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_725, data_out=>output_MAC_4_725);
	MAC_4_726: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_726, data_out=>output_MAC_4_726);
	MAC_4_727: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_727, data_out=>output_MAC_4_727);
	MAC_4_728: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_728, data_out=>output_MAC_4_728);
	MAC_4_729: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_729, data_out=>output_MAC_4_729);
	MAC_4_730: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_730, data_out=>output_MAC_4_730);
	MAC_4_731: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_731, data_out=>output_MAC_4_731);
	MAC_4_732: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_732, data_out=>output_MAC_4_732);
	MAC_4_733: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_733, data_out=>output_MAC_4_733);
	MAC_4_734: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_734, data_out=>output_MAC_4_734);
	MAC_4_735: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_735, data_out=>output_MAC_4_735);
	MAC_4_736: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_736, data_out=>output_MAC_4_736);
	MAC_4_737: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_737, data_out=>output_MAC_4_737);
	MAC_4_738: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_738, data_out=>output_MAC_4_738);
	MAC_4_739: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_739, data_out=>output_MAC_4_739);
	MAC_4_740: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_740, data_out=>output_MAC_4_740);
	MAC_4_741: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_741, data_out=>output_MAC_4_741);
	MAC_4_742: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_742, data_out=>output_MAC_4_742);
	MAC_4_743: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_743, data_out=>output_MAC_4_743);
	MAC_4_744: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_744, data_out=>output_MAC_4_744);
	MAC_4_745: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_745, data_out=>output_MAC_4_745);
	MAC_4_746: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_746, data_out=>output_MAC_4_746);
	MAC_4_747: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_747, data_out=>output_MAC_4_747);
	MAC_4_748: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_748, data_out=>output_MAC_4_748);
	MAC_4_749: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_749, data_out=>output_MAC_4_749);
	MAC_4_750: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_750, data_out=>output_MAC_4_750);
	MAC_4_751: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_751, data_out=>output_MAC_4_751);
	MAC_4_752: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_752, data_out=>output_MAC_4_752);
	MAC_4_753: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_753, data_out=>output_MAC_4_753);
	MAC_4_754: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_754, data_out=>output_MAC_4_754);
	MAC_4_755: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_755, data_out=>output_MAC_4_755);
	MAC_4_756: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_756, data_out=>output_MAC_4_756);
	MAC_4_757: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_757, data_out=>output_MAC_4_757);
	MAC_4_758: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_758, data_out=>output_MAC_4_758);
	MAC_4_759: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_759, data_out=>output_MAC_4_759);
	MAC_4_760: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_760, data_out=>output_MAC_4_760);
	MAC_4_761: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_761, data_out=>output_MAC_4_761);
	MAC_4_762: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_762, data_out=>output_MAC_4_762);
	MAC_4_763: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_763, data_out=>output_MAC_4_763);
	MAC_4_764: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_764, data_out=>output_MAC_4_764);
	MAC_4_765: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_765, data_out=>output_MAC_4_765);
	MAC_4_766: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_766, data_out=>output_MAC_4_766);
	MAC_4_767: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_4, data_in_B=>input_col_767, data_out=>output_MAC_4_767);
	MAC_5_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_0, data_out=>output_MAC_5_0);
	MAC_5_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_1, data_out=>output_MAC_5_1);
	MAC_5_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_2, data_out=>output_MAC_5_2);
	MAC_5_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_3, data_out=>output_MAC_5_3);
	MAC_5_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_4, data_out=>output_MAC_5_4);
	MAC_5_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_5, data_out=>output_MAC_5_5);
	MAC_5_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_6, data_out=>output_MAC_5_6);
	MAC_5_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_7, data_out=>output_MAC_5_7);
	MAC_5_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_8, data_out=>output_MAC_5_8);
	MAC_5_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_9, data_out=>output_MAC_5_9);
	MAC_5_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_10, data_out=>output_MAC_5_10);
	MAC_5_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_11, data_out=>output_MAC_5_11);
	MAC_5_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_12, data_out=>output_MAC_5_12);
	MAC_5_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_13, data_out=>output_MAC_5_13);
	MAC_5_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_14, data_out=>output_MAC_5_14);
	MAC_5_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_15, data_out=>output_MAC_5_15);
	MAC_5_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_16, data_out=>output_MAC_5_16);
	MAC_5_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_17, data_out=>output_MAC_5_17);
	MAC_5_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_18, data_out=>output_MAC_5_18);
	MAC_5_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_19, data_out=>output_MAC_5_19);
	MAC_5_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_20, data_out=>output_MAC_5_20);
	MAC_5_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_21, data_out=>output_MAC_5_21);
	MAC_5_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_22, data_out=>output_MAC_5_22);
	MAC_5_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_23, data_out=>output_MAC_5_23);
	MAC_5_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_24, data_out=>output_MAC_5_24);
	MAC_5_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_25, data_out=>output_MAC_5_25);
	MAC_5_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_26, data_out=>output_MAC_5_26);
	MAC_5_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_27, data_out=>output_MAC_5_27);
	MAC_5_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_28, data_out=>output_MAC_5_28);
	MAC_5_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_29, data_out=>output_MAC_5_29);
	MAC_5_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_30, data_out=>output_MAC_5_30);
	MAC_5_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_31, data_out=>output_MAC_5_31);
	MAC_5_32: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_32, data_out=>output_MAC_5_32);
	MAC_5_33: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_33, data_out=>output_MAC_5_33);
	MAC_5_34: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_34, data_out=>output_MAC_5_34);
	MAC_5_35: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_35, data_out=>output_MAC_5_35);
	MAC_5_36: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_36, data_out=>output_MAC_5_36);
	MAC_5_37: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_37, data_out=>output_MAC_5_37);
	MAC_5_38: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_38, data_out=>output_MAC_5_38);
	MAC_5_39: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_39, data_out=>output_MAC_5_39);
	MAC_5_40: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_40, data_out=>output_MAC_5_40);
	MAC_5_41: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_41, data_out=>output_MAC_5_41);
	MAC_5_42: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_42, data_out=>output_MAC_5_42);
	MAC_5_43: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_43, data_out=>output_MAC_5_43);
	MAC_5_44: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_44, data_out=>output_MAC_5_44);
	MAC_5_45: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_45, data_out=>output_MAC_5_45);
	MAC_5_46: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_46, data_out=>output_MAC_5_46);
	MAC_5_47: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_47, data_out=>output_MAC_5_47);
	MAC_5_48: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_48, data_out=>output_MAC_5_48);
	MAC_5_49: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_49, data_out=>output_MAC_5_49);
	MAC_5_50: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_50, data_out=>output_MAC_5_50);
	MAC_5_51: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_51, data_out=>output_MAC_5_51);
	MAC_5_52: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_52, data_out=>output_MAC_5_52);
	MAC_5_53: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_53, data_out=>output_MAC_5_53);
	MAC_5_54: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_54, data_out=>output_MAC_5_54);
	MAC_5_55: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_55, data_out=>output_MAC_5_55);
	MAC_5_56: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_56, data_out=>output_MAC_5_56);
	MAC_5_57: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_57, data_out=>output_MAC_5_57);
	MAC_5_58: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_58, data_out=>output_MAC_5_58);
	MAC_5_59: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_59, data_out=>output_MAC_5_59);
	MAC_5_60: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_60, data_out=>output_MAC_5_60);
	MAC_5_61: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_61, data_out=>output_MAC_5_61);
	MAC_5_62: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_62, data_out=>output_MAC_5_62);
	MAC_5_63: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_63, data_out=>output_MAC_5_63);
	MAC_5_64: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_64, data_out=>output_MAC_5_64);
	MAC_5_65: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_65, data_out=>output_MAC_5_65);
	MAC_5_66: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_66, data_out=>output_MAC_5_66);
	MAC_5_67: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_67, data_out=>output_MAC_5_67);
	MAC_5_68: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_68, data_out=>output_MAC_5_68);
	MAC_5_69: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_69, data_out=>output_MAC_5_69);
	MAC_5_70: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_70, data_out=>output_MAC_5_70);
	MAC_5_71: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_71, data_out=>output_MAC_5_71);
	MAC_5_72: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_72, data_out=>output_MAC_5_72);
	MAC_5_73: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_73, data_out=>output_MAC_5_73);
	MAC_5_74: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_74, data_out=>output_MAC_5_74);
	MAC_5_75: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_75, data_out=>output_MAC_5_75);
	MAC_5_76: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_76, data_out=>output_MAC_5_76);
	MAC_5_77: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_77, data_out=>output_MAC_5_77);
	MAC_5_78: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_78, data_out=>output_MAC_5_78);
	MAC_5_79: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_79, data_out=>output_MAC_5_79);
	MAC_5_80: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_80, data_out=>output_MAC_5_80);
	MAC_5_81: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_81, data_out=>output_MAC_5_81);
	MAC_5_82: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_82, data_out=>output_MAC_5_82);
	MAC_5_83: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_83, data_out=>output_MAC_5_83);
	MAC_5_84: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_84, data_out=>output_MAC_5_84);
	MAC_5_85: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_85, data_out=>output_MAC_5_85);
	MAC_5_86: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_86, data_out=>output_MAC_5_86);
	MAC_5_87: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_87, data_out=>output_MAC_5_87);
	MAC_5_88: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_88, data_out=>output_MAC_5_88);
	MAC_5_89: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_89, data_out=>output_MAC_5_89);
	MAC_5_90: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_90, data_out=>output_MAC_5_90);
	MAC_5_91: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_91, data_out=>output_MAC_5_91);
	MAC_5_92: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_92, data_out=>output_MAC_5_92);
	MAC_5_93: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_93, data_out=>output_MAC_5_93);
	MAC_5_94: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_94, data_out=>output_MAC_5_94);
	MAC_5_95: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_95, data_out=>output_MAC_5_95);
	MAC_5_96: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_96, data_out=>output_MAC_5_96);
	MAC_5_97: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_97, data_out=>output_MAC_5_97);
	MAC_5_98: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_98, data_out=>output_MAC_5_98);
	MAC_5_99: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_99, data_out=>output_MAC_5_99);
	MAC_5_100: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_100, data_out=>output_MAC_5_100);
	MAC_5_101: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_101, data_out=>output_MAC_5_101);
	MAC_5_102: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_102, data_out=>output_MAC_5_102);
	MAC_5_103: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_103, data_out=>output_MAC_5_103);
	MAC_5_104: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_104, data_out=>output_MAC_5_104);
	MAC_5_105: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_105, data_out=>output_MAC_5_105);
	MAC_5_106: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_106, data_out=>output_MAC_5_106);
	MAC_5_107: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_107, data_out=>output_MAC_5_107);
	MAC_5_108: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_108, data_out=>output_MAC_5_108);
	MAC_5_109: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_109, data_out=>output_MAC_5_109);
	MAC_5_110: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_110, data_out=>output_MAC_5_110);
	MAC_5_111: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_111, data_out=>output_MAC_5_111);
	MAC_5_112: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_112, data_out=>output_MAC_5_112);
	MAC_5_113: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_113, data_out=>output_MAC_5_113);
	MAC_5_114: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_114, data_out=>output_MAC_5_114);
	MAC_5_115: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_115, data_out=>output_MAC_5_115);
	MAC_5_116: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_116, data_out=>output_MAC_5_116);
	MAC_5_117: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_117, data_out=>output_MAC_5_117);
	MAC_5_118: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_118, data_out=>output_MAC_5_118);
	MAC_5_119: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_119, data_out=>output_MAC_5_119);
	MAC_5_120: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_120, data_out=>output_MAC_5_120);
	MAC_5_121: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_121, data_out=>output_MAC_5_121);
	MAC_5_122: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_122, data_out=>output_MAC_5_122);
	MAC_5_123: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_123, data_out=>output_MAC_5_123);
	MAC_5_124: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_124, data_out=>output_MAC_5_124);
	MAC_5_125: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_125, data_out=>output_MAC_5_125);
	MAC_5_126: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_126, data_out=>output_MAC_5_126);
	MAC_5_127: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_127, data_out=>output_MAC_5_127);
	MAC_5_128: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_128, data_out=>output_MAC_5_128);
	MAC_5_129: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_129, data_out=>output_MAC_5_129);
	MAC_5_130: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_130, data_out=>output_MAC_5_130);
	MAC_5_131: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_131, data_out=>output_MAC_5_131);
	MAC_5_132: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_132, data_out=>output_MAC_5_132);
	MAC_5_133: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_133, data_out=>output_MAC_5_133);
	MAC_5_134: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_134, data_out=>output_MAC_5_134);
	MAC_5_135: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_135, data_out=>output_MAC_5_135);
	MAC_5_136: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_136, data_out=>output_MAC_5_136);
	MAC_5_137: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_137, data_out=>output_MAC_5_137);
	MAC_5_138: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_138, data_out=>output_MAC_5_138);
	MAC_5_139: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_139, data_out=>output_MAC_5_139);
	MAC_5_140: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_140, data_out=>output_MAC_5_140);
	MAC_5_141: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_141, data_out=>output_MAC_5_141);
	MAC_5_142: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_142, data_out=>output_MAC_5_142);
	MAC_5_143: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_143, data_out=>output_MAC_5_143);
	MAC_5_144: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_144, data_out=>output_MAC_5_144);
	MAC_5_145: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_145, data_out=>output_MAC_5_145);
	MAC_5_146: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_146, data_out=>output_MAC_5_146);
	MAC_5_147: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_147, data_out=>output_MAC_5_147);
	MAC_5_148: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_148, data_out=>output_MAC_5_148);
	MAC_5_149: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_149, data_out=>output_MAC_5_149);
	MAC_5_150: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_150, data_out=>output_MAC_5_150);
	MAC_5_151: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_151, data_out=>output_MAC_5_151);
	MAC_5_152: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_152, data_out=>output_MAC_5_152);
	MAC_5_153: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_153, data_out=>output_MAC_5_153);
	MAC_5_154: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_154, data_out=>output_MAC_5_154);
	MAC_5_155: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_155, data_out=>output_MAC_5_155);
	MAC_5_156: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_156, data_out=>output_MAC_5_156);
	MAC_5_157: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_157, data_out=>output_MAC_5_157);
	MAC_5_158: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_158, data_out=>output_MAC_5_158);
	MAC_5_159: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_159, data_out=>output_MAC_5_159);
	MAC_5_160: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_160, data_out=>output_MAC_5_160);
	MAC_5_161: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_161, data_out=>output_MAC_5_161);
	MAC_5_162: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_162, data_out=>output_MAC_5_162);
	MAC_5_163: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_163, data_out=>output_MAC_5_163);
	MAC_5_164: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_164, data_out=>output_MAC_5_164);
	MAC_5_165: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_165, data_out=>output_MAC_5_165);
	MAC_5_166: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_166, data_out=>output_MAC_5_166);
	MAC_5_167: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_167, data_out=>output_MAC_5_167);
	MAC_5_168: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_168, data_out=>output_MAC_5_168);
	MAC_5_169: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_169, data_out=>output_MAC_5_169);
	MAC_5_170: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_170, data_out=>output_MAC_5_170);
	MAC_5_171: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_171, data_out=>output_MAC_5_171);
	MAC_5_172: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_172, data_out=>output_MAC_5_172);
	MAC_5_173: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_173, data_out=>output_MAC_5_173);
	MAC_5_174: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_174, data_out=>output_MAC_5_174);
	MAC_5_175: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_175, data_out=>output_MAC_5_175);
	MAC_5_176: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_176, data_out=>output_MAC_5_176);
	MAC_5_177: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_177, data_out=>output_MAC_5_177);
	MAC_5_178: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_178, data_out=>output_MAC_5_178);
	MAC_5_179: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_179, data_out=>output_MAC_5_179);
	MAC_5_180: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_180, data_out=>output_MAC_5_180);
	MAC_5_181: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_181, data_out=>output_MAC_5_181);
	MAC_5_182: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_182, data_out=>output_MAC_5_182);
	MAC_5_183: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_183, data_out=>output_MAC_5_183);
	MAC_5_184: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_184, data_out=>output_MAC_5_184);
	MAC_5_185: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_185, data_out=>output_MAC_5_185);
	MAC_5_186: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_186, data_out=>output_MAC_5_186);
	MAC_5_187: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_187, data_out=>output_MAC_5_187);
	MAC_5_188: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_188, data_out=>output_MAC_5_188);
	MAC_5_189: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_189, data_out=>output_MAC_5_189);
	MAC_5_190: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_190, data_out=>output_MAC_5_190);
	MAC_5_191: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_191, data_out=>output_MAC_5_191);
	MAC_5_192: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_192, data_out=>output_MAC_5_192);
	MAC_5_193: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_193, data_out=>output_MAC_5_193);
	MAC_5_194: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_194, data_out=>output_MAC_5_194);
	MAC_5_195: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_195, data_out=>output_MAC_5_195);
	MAC_5_196: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_196, data_out=>output_MAC_5_196);
	MAC_5_197: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_197, data_out=>output_MAC_5_197);
	MAC_5_198: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_198, data_out=>output_MAC_5_198);
	MAC_5_199: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_199, data_out=>output_MAC_5_199);
	MAC_5_200: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_200, data_out=>output_MAC_5_200);
	MAC_5_201: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_201, data_out=>output_MAC_5_201);
	MAC_5_202: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_202, data_out=>output_MAC_5_202);
	MAC_5_203: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_203, data_out=>output_MAC_5_203);
	MAC_5_204: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_204, data_out=>output_MAC_5_204);
	MAC_5_205: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_205, data_out=>output_MAC_5_205);
	MAC_5_206: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_206, data_out=>output_MAC_5_206);
	MAC_5_207: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_207, data_out=>output_MAC_5_207);
	MAC_5_208: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_208, data_out=>output_MAC_5_208);
	MAC_5_209: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_209, data_out=>output_MAC_5_209);
	MAC_5_210: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_210, data_out=>output_MAC_5_210);
	MAC_5_211: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_211, data_out=>output_MAC_5_211);
	MAC_5_212: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_212, data_out=>output_MAC_5_212);
	MAC_5_213: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_213, data_out=>output_MAC_5_213);
	MAC_5_214: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_214, data_out=>output_MAC_5_214);
	MAC_5_215: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_215, data_out=>output_MAC_5_215);
	MAC_5_216: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_216, data_out=>output_MAC_5_216);
	MAC_5_217: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_217, data_out=>output_MAC_5_217);
	MAC_5_218: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_218, data_out=>output_MAC_5_218);
	MAC_5_219: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_219, data_out=>output_MAC_5_219);
	MAC_5_220: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_220, data_out=>output_MAC_5_220);
	MAC_5_221: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_221, data_out=>output_MAC_5_221);
	MAC_5_222: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_222, data_out=>output_MAC_5_222);
	MAC_5_223: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_223, data_out=>output_MAC_5_223);
	MAC_5_224: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_224, data_out=>output_MAC_5_224);
	MAC_5_225: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_225, data_out=>output_MAC_5_225);
	MAC_5_226: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_226, data_out=>output_MAC_5_226);
	MAC_5_227: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_227, data_out=>output_MAC_5_227);
	MAC_5_228: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_228, data_out=>output_MAC_5_228);
	MAC_5_229: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_229, data_out=>output_MAC_5_229);
	MAC_5_230: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_230, data_out=>output_MAC_5_230);
	MAC_5_231: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_231, data_out=>output_MAC_5_231);
	MAC_5_232: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_232, data_out=>output_MAC_5_232);
	MAC_5_233: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_233, data_out=>output_MAC_5_233);
	MAC_5_234: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_234, data_out=>output_MAC_5_234);
	MAC_5_235: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_235, data_out=>output_MAC_5_235);
	MAC_5_236: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_236, data_out=>output_MAC_5_236);
	MAC_5_237: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_237, data_out=>output_MAC_5_237);
	MAC_5_238: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_238, data_out=>output_MAC_5_238);
	MAC_5_239: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_239, data_out=>output_MAC_5_239);
	MAC_5_240: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_240, data_out=>output_MAC_5_240);
	MAC_5_241: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_241, data_out=>output_MAC_5_241);
	MAC_5_242: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_242, data_out=>output_MAC_5_242);
	MAC_5_243: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_243, data_out=>output_MAC_5_243);
	MAC_5_244: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_244, data_out=>output_MAC_5_244);
	MAC_5_245: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_245, data_out=>output_MAC_5_245);
	MAC_5_246: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_246, data_out=>output_MAC_5_246);
	MAC_5_247: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_247, data_out=>output_MAC_5_247);
	MAC_5_248: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_248, data_out=>output_MAC_5_248);
	MAC_5_249: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_249, data_out=>output_MAC_5_249);
	MAC_5_250: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_250, data_out=>output_MAC_5_250);
	MAC_5_251: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_251, data_out=>output_MAC_5_251);
	MAC_5_252: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_252, data_out=>output_MAC_5_252);
	MAC_5_253: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_253, data_out=>output_MAC_5_253);
	MAC_5_254: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_254, data_out=>output_MAC_5_254);
	MAC_5_255: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_255, data_out=>output_MAC_5_255);
	MAC_5_256: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_256, data_out=>output_MAC_5_256);
	MAC_5_257: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_257, data_out=>output_MAC_5_257);
	MAC_5_258: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_258, data_out=>output_MAC_5_258);
	MAC_5_259: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_259, data_out=>output_MAC_5_259);
	MAC_5_260: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_260, data_out=>output_MAC_5_260);
	MAC_5_261: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_261, data_out=>output_MAC_5_261);
	MAC_5_262: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_262, data_out=>output_MAC_5_262);
	MAC_5_263: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_263, data_out=>output_MAC_5_263);
	MAC_5_264: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_264, data_out=>output_MAC_5_264);
	MAC_5_265: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_265, data_out=>output_MAC_5_265);
	MAC_5_266: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_266, data_out=>output_MAC_5_266);
	MAC_5_267: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_267, data_out=>output_MAC_5_267);
	MAC_5_268: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_268, data_out=>output_MAC_5_268);
	MAC_5_269: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_269, data_out=>output_MAC_5_269);
	MAC_5_270: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_270, data_out=>output_MAC_5_270);
	MAC_5_271: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_271, data_out=>output_MAC_5_271);
	MAC_5_272: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_272, data_out=>output_MAC_5_272);
	MAC_5_273: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_273, data_out=>output_MAC_5_273);
	MAC_5_274: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_274, data_out=>output_MAC_5_274);
	MAC_5_275: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_275, data_out=>output_MAC_5_275);
	MAC_5_276: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_276, data_out=>output_MAC_5_276);
	MAC_5_277: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_277, data_out=>output_MAC_5_277);
	MAC_5_278: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_278, data_out=>output_MAC_5_278);
	MAC_5_279: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_279, data_out=>output_MAC_5_279);
	MAC_5_280: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_280, data_out=>output_MAC_5_280);
	MAC_5_281: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_281, data_out=>output_MAC_5_281);
	MAC_5_282: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_282, data_out=>output_MAC_5_282);
	MAC_5_283: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_283, data_out=>output_MAC_5_283);
	MAC_5_284: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_284, data_out=>output_MAC_5_284);
	MAC_5_285: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_285, data_out=>output_MAC_5_285);
	MAC_5_286: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_286, data_out=>output_MAC_5_286);
	MAC_5_287: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_287, data_out=>output_MAC_5_287);
	MAC_5_288: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_288, data_out=>output_MAC_5_288);
	MAC_5_289: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_289, data_out=>output_MAC_5_289);
	MAC_5_290: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_290, data_out=>output_MAC_5_290);
	MAC_5_291: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_291, data_out=>output_MAC_5_291);
	MAC_5_292: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_292, data_out=>output_MAC_5_292);
	MAC_5_293: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_293, data_out=>output_MAC_5_293);
	MAC_5_294: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_294, data_out=>output_MAC_5_294);
	MAC_5_295: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_295, data_out=>output_MAC_5_295);
	MAC_5_296: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_296, data_out=>output_MAC_5_296);
	MAC_5_297: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_297, data_out=>output_MAC_5_297);
	MAC_5_298: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_298, data_out=>output_MAC_5_298);
	MAC_5_299: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_299, data_out=>output_MAC_5_299);
	MAC_5_300: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_300, data_out=>output_MAC_5_300);
	MAC_5_301: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_301, data_out=>output_MAC_5_301);
	MAC_5_302: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_302, data_out=>output_MAC_5_302);
	MAC_5_303: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_303, data_out=>output_MAC_5_303);
	MAC_5_304: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_304, data_out=>output_MAC_5_304);
	MAC_5_305: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_305, data_out=>output_MAC_5_305);
	MAC_5_306: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_306, data_out=>output_MAC_5_306);
	MAC_5_307: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_307, data_out=>output_MAC_5_307);
	MAC_5_308: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_308, data_out=>output_MAC_5_308);
	MAC_5_309: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_309, data_out=>output_MAC_5_309);
	MAC_5_310: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_310, data_out=>output_MAC_5_310);
	MAC_5_311: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_311, data_out=>output_MAC_5_311);
	MAC_5_312: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_312, data_out=>output_MAC_5_312);
	MAC_5_313: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_313, data_out=>output_MAC_5_313);
	MAC_5_314: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_314, data_out=>output_MAC_5_314);
	MAC_5_315: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_315, data_out=>output_MAC_5_315);
	MAC_5_316: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_316, data_out=>output_MAC_5_316);
	MAC_5_317: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_317, data_out=>output_MAC_5_317);
	MAC_5_318: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_318, data_out=>output_MAC_5_318);
	MAC_5_319: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_319, data_out=>output_MAC_5_319);
	MAC_5_320: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_320, data_out=>output_MAC_5_320);
	MAC_5_321: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_321, data_out=>output_MAC_5_321);
	MAC_5_322: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_322, data_out=>output_MAC_5_322);
	MAC_5_323: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_323, data_out=>output_MAC_5_323);
	MAC_5_324: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_324, data_out=>output_MAC_5_324);
	MAC_5_325: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_325, data_out=>output_MAC_5_325);
	MAC_5_326: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_326, data_out=>output_MAC_5_326);
	MAC_5_327: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_327, data_out=>output_MAC_5_327);
	MAC_5_328: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_328, data_out=>output_MAC_5_328);
	MAC_5_329: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_329, data_out=>output_MAC_5_329);
	MAC_5_330: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_330, data_out=>output_MAC_5_330);
	MAC_5_331: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_331, data_out=>output_MAC_5_331);
	MAC_5_332: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_332, data_out=>output_MAC_5_332);
	MAC_5_333: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_333, data_out=>output_MAC_5_333);
	MAC_5_334: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_334, data_out=>output_MAC_5_334);
	MAC_5_335: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_335, data_out=>output_MAC_5_335);
	MAC_5_336: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_336, data_out=>output_MAC_5_336);
	MAC_5_337: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_337, data_out=>output_MAC_5_337);
	MAC_5_338: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_338, data_out=>output_MAC_5_338);
	MAC_5_339: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_339, data_out=>output_MAC_5_339);
	MAC_5_340: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_340, data_out=>output_MAC_5_340);
	MAC_5_341: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_341, data_out=>output_MAC_5_341);
	MAC_5_342: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_342, data_out=>output_MAC_5_342);
	MAC_5_343: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_343, data_out=>output_MAC_5_343);
	MAC_5_344: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_344, data_out=>output_MAC_5_344);
	MAC_5_345: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_345, data_out=>output_MAC_5_345);
	MAC_5_346: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_346, data_out=>output_MAC_5_346);
	MAC_5_347: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_347, data_out=>output_MAC_5_347);
	MAC_5_348: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_348, data_out=>output_MAC_5_348);
	MAC_5_349: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_349, data_out=>output_MAC_5_349);
	MAC_5_350: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_350, data_out=>output_MAC_5_350);
	MAC_5_351: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_351, data_out=>output_MAC_5_351);
	MAC_5_352: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_352, data_out=>output_MAC_5_352);
	MAC_5_353: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_353, data_out=>output_MAC_5_353);
	MAC_5_354: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_354, data_out=>output_MAC_5_354);
	MAC_5_355: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_355, data_out=>output_MAC_5_355);
	MAC_5_356: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_356, data_out=>output_MAC_5_356);
	MAC_5_357: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_357, data_out=>output_MAC_5_357);
	MAC_5_358: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_358, data_out=>output_MAC_5_358);
	MAC_5_359: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_359, data_out=>output_MAC_5_359);
	MAC_5_360: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_360, data_out=>output_MAC_5_360);
	MAC_5_361: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_361, data_out=>output_MAC_5_361);
	MAC_5_362: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_362, data_out=>output_MAC_5_362);
	MAC_5_363: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_363, data_out=>output_MAC_5_363);
	MAC_5_364: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_364, data_out=>output_MAC_5_364);
	MAC_5_365: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_365, data_out=>output_MAC_5_365);
	MAC_5_366: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_366, data_out=>output_MAC_5_366);
	MAC_5_367: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_367, data_out=>output_MAC_5_367);
	MAC_5_368: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_368, data_out=>output_MAC_5_368);
	MAC_5_369: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_369, data_out=>output_MAC_5_369);
	MAC_5_370: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_370, data_out=>output_MAC_5_370);
	MAC_5_371: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_371, data_out=>output_MAC_5_371);
	MAC_5_372: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_372, data_out=>output_MAC_5_372);
	MAC_5_373: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_373, data_out=>output_MAC_5_373);
	MAC_5_374: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_374, data_out=>output_MAC_5_374);
	MAC_5_375: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_375, data_out=>output_MAC_5_375);
	MAC_5_376: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_376, data_out=>output_MAC_5_376);
	MAC_5_377: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_377, data_out=>output_MAC_5_377);
	MAC_5_378: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_378, data_out=>output_MAC_5_378);
	MAC_5_379: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_379, data_out=>output_MAC_5_379);
	MAC_5_380: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_380, data_out=>output_MAC_5_380);
	MAC_5_381: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_381, data_out=>output_MAC_5_381);
	MAC_5_382: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_382, data_out=>output_MAC_5_382);
	MAC_5_383: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_383, data_out=>output_MAC_5_383);
	MAC_5_384: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_384, data_out=>output_MAC_5_384);
	MAC_5_385: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_385, data_out=>output_MAC_5_385);
	MAC_5_386: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_386, data_out=>output_MAC_5_386);
	MAC_5_387: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_387, data_out=>output_MAC_5_387);
	MAC_5_388: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_388, data_out=>output_MAC_5_388);
	MAC_5_389: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_389, data_out=>output_MAC_5_389);
	MAC_5_390: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_390, data_out=>output_MAC_5_390);
	MAC_5_391: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_391, data_out=>output_MAC_5_391);
	MAC_5_392: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_392, data_out=>output_MAC_5_392);
	MAC_5_393: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_393, data_out=>output_MAC_5_393);
	MAC_5_394: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_394, data_out=>output_MAC_5_394);
	MAC_5_395: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_395, data_out=>output_MAC_5_395);
	MAC_5_396: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_396, data_out=>output_MAC_5_396);
	MAC_5_397: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_397, data_out=>output_MAC_5_397);
	MAC_5_398: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_398, data_out=>output_MAC_5_398);
	MAC_5_399: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_399, data_out=>output_MAC_5_399);
	MAC_5_400: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_400, data_out=>output_MAC_5_400);
	MAC_5_401: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_401, data_out=>output_MAC_5_401);
	MAC_5_402: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_402, data_out=>output_MAC_5_402);
	MAC_5_403: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_403, data_out=>output_MAC_5_403);
	MAC_5_404: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_404, data_out=>output_MAC_5_404);
	MAC_5_405: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_405, data_out=>output_MAC_5_405);
	MAC_5_406: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_406, data_out=>output_MAC_5_406);
	MAC_5_407: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_407, data_out=>output_MAC_5_407);
	MAC_5_408: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_408, data_out=>output_MAC_5_408);
	MAC_5_409: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_409, data_out=>output_MAC_5_409);
	MAC_5_410: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_410, data_out=>output_MAC_5_410);
	MAC_5_411: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_411, data_out=>output_MAC_5_411);
	MAC_5_412: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_412, data_out=>output_MAC_5_412);
	MAC_5_413: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_413, data_out=>output_MAC_5_413);
	MAC_5_414: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_414, data_out=>output_MAC_5_414);
	MAC_5_415: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_415, data_out=>output_MAC_5_415);
	MAC_5_416: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_416, data_out=>output_MAC_5_416);
	MAC_5_417: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_417, data_out=>output_MAC_5_417);
	MAC_5_418: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_418, data_out=>output_MAC_5_418);
	MAC_5_419: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_419, data_out=>output_MAC_5_419);
	MAC_5_420: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_420, data_out=>output_MAC_5_420);
	MAC_5_421: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_421, data_out=>output_MAC_5_421);
	MAC_5_422: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_422, data_out=>output_MAC_5_422);
	MAC_5_423: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_423, data_out=>output_MAC_5_423);
	MAC_5_424: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_424, data_out=>output_MAC_5_424);
	MAC_5_425: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_425, data_out=>output_MAC_5_425);
	MAC_5_426: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_426, data_out=>output_MAC_5_426);
	MAC_5_427: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_427, data_out=>output_MAC_5_427);
	MAC_5_428: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_428, data_out=>output_MAC_5_428);
	MAC_5_429: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_429, data_out=>output_MAC_5_429);
	MAC_5_430: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_430, data_out=>output_MAC_5_430);
	MAC_5_431: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_431, data_out=>output_MAC_5_431);
	MAC_5_432: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_432, data_out=>output_MAC_5_432);
	MAC_5_433: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_433, data_out=>output_MAC_5_433);
	MAC_5_434: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_434, data_out=>output_MAC_5_434);
	MAC_5_435: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_435, data_out=>output_MAC_5_435);
	MAC_5_436: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_436, data_out=>output_MAC_5_436);
	MAC_5_437: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_437, data_out=>output_MAC_5_437);
	MAC_5_438: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_438, data_out=>output_MAC_5_438);
	MAC_5_439: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_439, data_out=>output_MAC_5_439);
	MAC_5_440: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_440, data_out=>output_MAC_5_440);
	MAC_5_441: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_441, data_out=>output_MAC_5_441);
	MAC_5_442: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_442, data_out=>output_MAC_5_442);
	MAC_5_443: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_443, data_out=>output_MAC_5_443);
	MAC_5_444: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_444, data_out=>output_MAC_5_444);
	MAC_5_445: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_445, data_out=>output_MAC_5_445);
	MAC_5_446: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_446, data_out=>output_MAC_5_446);
	MAC_5_447: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_447, data_out=>output_MAC_5_447);
	MAC_5_448: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_448, data_out=>output_MAC_5_448);
	MAC_5_449: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_449, data_out=>output_MAC_5_449);
	MAC_5_450: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_450, data_out=>output_MAC_5_450);
	MAC_5_451: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_451, data_out=>output_MAC_5_451);
	MAC_5_452: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_452, data_out=>output_MAC_5_452);
	MAC_5_453: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_453, data_out=>output_MAC_5_453);
	MAC_5_454: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_454, data_out=>output_MAC_5_454);
	MAC_5_455: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_455, data_out=>output_MAC_5_455);
	MAC_5_456: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_456, data_out=>output_MAC_5_456);
	MAC_5_457: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_457, data_out=>output_MAC_5_457);
	MAC_5_458: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_458, data_out=>output_MAC_5_458);
	MAC_5_459: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_459, data_out=>output_MAC_5_459);
	MAC_5_460: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_460, data_out=>output_MAC_5_460);
	MAC_5_461: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_461, data_out=>output_MAC_5_461);
	MAC_5_462: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_462, data_out=>output_MAC_5_462);
	MAC_5_463: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_463, data_out=>output_MAC_5_463);
	MAC_5_464: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_464, data_out=>output_MAC_5_464);
	MAC_5_465: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_465, data_out=>output_MAC_5_465);
	MAC_5_466: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_466, data_out=>output_MAC_5_466);
	MAC_5_467: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_467, data_out=>output_MAC_5_467);
	MAC_5_468: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_468, data_out=>output_MAC_5_468);
	MAC_5_469: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_469, data_out=>output_MAC_5_469);
	MAC_5_470: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_470, data_out=>output_MAC_5_470);
	MAC_5_471: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_471, data_out=>output_MAC_5_471);
	MAC_5_472: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_472, data_out=>output_MAC_5_472);
	MAC_5_473: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_473, data_out=>output_MAC_5_473);
	MAC_5_474: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_474, data_out=>output_MAC_5_474);
	MAC_5_475: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_475, data_out=>output_MAC_5_475);
	MAC_5_476: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_476, data_out=>output_MAC_5_476);
	MAC_5_477: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_477, data_out=>output_MAC_5_477);
	MAC_5_478: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_478, data_out=>output_MAC_5_478);
	MAC_5_479: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_479, data_out=>output_MAC_5_479);
	MAC_5_480: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_480, data_out=>output_MAC_5_480);
	MAC_5_481: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_481, data_out=>output_MAC_5_481);
	MAC_5_482: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_482, data_out=>output_MAC_5_482);
	MAC_5_483: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_483, data_out=>output_MAC_5_483);
	MAC_5_484: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_484, data_out=>output_MAC_5_484);
	MAC_5_485: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_485, data_out=>output_MAC_5_485);
	MAC_5_486: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_486, data_out=>output_MAC_5_486);
	MAC_5_487: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_487, data_out=>output_MAC_5_487);
	MAC_5_488: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_488, data_out=>output_MAC_5_488);
	MAC_5_489: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_489, data_out=>output_MAC_5_489);
	MAC_5_490: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_490, data_out=>output_MAC_5_490);
	MAC_5_491: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_491, data_out=>output_MAC_5_491);
	MAC_5_492: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_492, data_out=>output_MAC_5_492);
	MAC_5_493: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_493, data_out=>output_MAC_5_493);
	MAC_5_494: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_494, data_out=>output_MAC_5_494);
	MAC_5_495: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_495, data_out=>output_MAC_5_495);
	MAC_5_496: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_496, data_out=>output_MAC_5_496);
	MAC_5_497: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_497, data_out=>output_MAC_5_497);
	MAC_5_498: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_498, data_out=>output_MAC_5_498);
	MAC_5_499: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_499, data_out=>output_MAC_5_499);
	MAC_5_500: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_500, data_out=>output_MAC_5_500);
	MAC_5_501: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_501, data_out=>output_MAC_5_501);
	MAC_5_502: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_502, data_out=>output_MAC_5_502);
	MAC_5_503: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_503, data_out=>output_MAC_5_503);
	MAC_5_504: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_504, data_out=>output_MAC_5_504);
	MAC_5_505: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_505, data_out=>output_MAC_5_505);
	MAC_5_506: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_506, data_out=>output_MAC_5_506);
	MAC_5_507: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_507, data_out=>output_MAC_5_507);
	MAC_5_508: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_508, data_out=>output_MAC_5_508);
	MAC_5_509: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_509, data_out=>output_MAC_5_509);
	MAC_5_510: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_510, data_out=>output_MAC_5_510);
	MAC_5_511: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_511, data_out=>output_MAC_5_511);
	MAC_5_512: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_512, data_out=>output_MAC_5_512);
	MAC_5_513: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_513, data_out=>output_MAC_5_513);
	MAC_5_514: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_514, data_out=>output_MAC_5_514);
	MAC_5_515: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_515, data_out=>output_MAC_5_515);
	MAC_5_516: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_516, data_out=>output_MAC_5_516);
	MAC_5_517: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_517, data_out=>output_MAC_5_517);
	MAC_5_518: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_518, data_out=>output_MAC_5_518);
	MAC_5_519: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_519, data_out=>output_MAC_5_519);
	MAC_5_520: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_520, data_out=>output_MAC_5_520);
	MAC_5_521: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_521, data_out=>output_MAC_5_521);
	MAC_5_522: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_522, data_out=>output_MAC_5_522);
	MAC_5_523: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_523, data_out=>output_MAC_5_523);
	MAC_5_524: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_524, data_out=>output_MAC_5_524);
	MAC_5_525: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_525, data_out=>output_MAC_5_525);
	MAC_5_526: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_526, data_out=>output_MAC_5_526);
	MAC_5_527: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_527, data_out=>output_MAC_5_527);
	MAC_5_528: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_528, data_out=>output_MAC_5_528);
	MAC_5_529: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_529, data_out=>output_MAC_5_529);
	MAC_5_530: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_530, data_out=>output_MAC_5_530);
	MAC_5_531: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_531, data_out=>output_MAC_5_531);
	MAC_5_532: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_532, data_out=>output_MAC_5_532);
	MAC_5_533: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_533, data_out=>output_MAC_5_533);
	MAC_5_534: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_534, data_out=>output_MAC_5_534);
	MAC_5_535: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_535, data_out=>output_MAC_5_535);
	MAC_5_536: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_536, data_out=>output_MAC_5_536);
	MAC_5_537: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_537, data_out=>output_MAC_5_537);
	MAC_5_538: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_538, data_out=>output_MAC_5_538);
	MAC_5_539: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_539, data_out=>output_MAC_5_539);
	MAC_5_540: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_540, data_out=>output_MAC_5_540);
	MAC_5_541: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_541, data_out=>output_MAC_5_541);
	MAC_5_542: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_542, data_out=>output_MAC_5_542);
	MAC_5_543: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_543, data_out=>output_MAC_5_543);
	MAC_5_544: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_544, data_out=>output_MAC_5_544);
	MAC_5_545: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_545, data_out=>output_MAC_5_545);
	MAC_5_546: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_546, data_out=>output_MAC_5_546);
	MAC_5_547: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_547, data_out=>output_MAC_5_547);
	MAC_5_548: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_548, data_out=>output_MAC_5_548);
	MAC_5_549: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_549, data_out=>output_MAC_5_549);
	MAC_5_550: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_550, data_out=>output_MAC_5_550);
	MAC_5_551: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_551, data_out=>output_MAC_5_551);
	MAC_5_552: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_552, data_out=>output_MAC_5_552);
	MAC_5_553: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_553, data_out=>output_MAC_5_553);
	MAC_5_554: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_554, data_out=>output_MAC_5_554);
	MAC_5_555: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_555, data_out=>output_MAC_5_555);
	MAC_5_556: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_556, data_out=>output_MAC_5_556);
	MAC_5_557: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_557, data_out=>output_MAC_5_557);
	MAC_5_558: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_558, data_out=>output_MAC_5_558);
	MAC_5_559: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_559, data_out=>output_MAC_5_559);
	MAC_5_560: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_560, data_out=>output_MAC_5_560);
	MAC_5_561: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_561, data_out=>output_MAC_5_561);
	MAC_5_562: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_562, data_out=>output_MAC_5_562);
	MAC_5_563: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_563, data_out=>output_MAC_5_563);
	MAC_5_564: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_564, data_out=>output_MAC_5_564);
	MAC_5_565: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_565, data_out=>output_MAC_5_565);
	MAC_5_566: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_566, data_out=>output_MAC_5_566);
	MAC_5_567: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_567, data_out=>output_MAC_5_567);
	MAC_5_568: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_568, data_out=>output_MAC_5_568);
	MAC_5_569: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_569, data_out=>output_MAC_5_569);
	MAC_5_570: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_570, data_out=>output_MAC_5_570);
	MAC_5_571: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_571, data_out=>output_MAC_5_571);
	MAC_5_572: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_572, data_out=>output_MAC_5_572);
	MAC_5_573: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_573, data_out=>output_MAC_5_573);
	MAC_5_574: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_574, data_out=>output_MAC_5_574);
	MAC_5_575: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_575, data_out=>output_MAC_5_575);
	MAC_5_576: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_576, data_out=>output_MAC_5_576);
	MAC_5_577: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_577, data_out=>output_MAC_5_577);
	MAC_5_578: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_578, data_out=>output_MAC_5_578);
	MAC_5_579: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_579, data_out=>output_MAC_5_579);
	MAC_5_580: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_580, data_out=>output_MAC_5_580);
	MAC_5_581: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_581, data_out=>output_MAC_5_581);
	MAC_5_582: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_582, data_out=>output_MAC_5_582);
	MAC_5_583: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_583, data_out=>output_MAC_5_583);
	MAC_5_584: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_584, data_out=>output_MAC_5_584);
	MAC_5_585: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_585, data_out=>output_MAC_5_585);
	MAC_5_586: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_586, data_out=>output_MAC_5_586);
	MAC_5_587: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_587, data_out=>output_MAC_5_587);
	MAC_5_588: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_588, data_out=>output_MAC_5_588);
	MAC_5_589: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_589, data_out=>output_MAC_5_589);
	MAC_5_590: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_590, data_out=>output_MAC_5_590);
	MAC_5_591: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_591, data_out=>output_MAC_5_591);
	MAC_5_592: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_592, data_out=>output_MAC_5_592);
	MAC_5_593: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_593, data_out=>output_MAC_5_593);
	MAC_5_594: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_594, data_out=>output_MAC_5_594);
	MAC_5_595: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_595, data_out=>output_MAC_5_595);
	MAC_5_596: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_596, data_out=>output_MAC_5_596);
	MAC_5_597: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_597, data_out=>output_MAC_5_597);
	MAC_5_598: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_598, data_out=>output_MAC_5_598);
	MAC_5_599: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_599, data_out=>output_MAC_5_599);
	MAC_5_600: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_600, data_out=>output_MAC_5_600);
	MAC_5_601: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_601, data_out=>output_MAC_5_601);
	MAC_5_602: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_602, data_out=>output_MAC_5_602);
	MAC_5_603: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_603, data_out=>output_MAC_5_603);
	MAC_5_604: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_604, data_out=>output_MAC_5_604);
	MAC_5_605: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_605, data_out=>output_MAC_5_605);
	MAC_5_606: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_606, data_out=>output_MAC_5_606);
	MAC_5_607: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_607, data_out=>output_MAC_5_607);
	MAC_5_608: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_608, data_out=>output_MAC_5_608);
	MAC_5_609: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_609, data_out=>output_MAC_5_609);
	MAC_5_610: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_610, data_out=>output_MAC_5_610);
	MAC_5_611: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_611, data_out=>output_MAC_5_611);
	MAC_5_612: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_612, data_out=>output_MAC_5_612);
	MAC_5_613: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_613, data_out=>output_MAC_5_613);
	MAC_5_614: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_614, data_out=>output_MAC_5_614);
	MAC_5_615: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_615, data_out=>output_MAC_5_615);
	MAC_5_616: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_616, data_out=>output_MAC_5_616);
	MAC_5_617: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_617, data_out=>output_MAC_5_617);
	MAC_5_618: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_618, data_out=>output_MAC_5_618);
	MAC_5_619: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_619, data_out=>output_MAC_5_619);
	MAC_5_620: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_620, data_out=>output_MAC_5_620);
	MAC_5_621: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_621, data_out=>output_MAC_5_621);
	MAC_5_622: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_622, data_out=>output_MAC_5_622);
	MAC_5_623: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_623, data_out=>output_MAC_5_623);
	MAC_5_624: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_624, data_out=>output_MAC_5_624);
	MAC_5_625: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_625, data_out=>output_MAC_5_625);
	MAC_5_626: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_626, data_out=>output_MAC_5_626);
	MAC_5_627: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_627, data_out=>output_MAC_5_627);
	MAC_5_628: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_628, data_out=>output_MAC_5_628);
	MAC_5_629: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_629, data_out=>output_MAC_5_629);
	MAC_5_630: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_630, data_out=>output_MAC_5_630);
	MAC_5_631: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_631, data_out=>output_MAC_5_631);
	MAC_5_632: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_632, data_out=>output_MAC_5_632);
	MAC_5_633: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_633, data_out=>output_MAC_5_633);
	MAC_5_634: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_634, data_out=>output_MAC_5_634);
	MAC_5_635: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_635, data_out=>output_MAC_5_635);
	MAC_5_636: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_636, data_out=>output_MAC_5_636);
	MAC_5_637: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_637, data_out=>output_MAC_5_637);
	MAC_5_638: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_638, data_out=>output_MAC_5_638);
	MAC_5_639: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_639, data_out=>output_MAC_5_639);
	MAC_5_640: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_640, data_out=>output_MAC_5_640);
	MAC_5_641: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_641, data_out=>output_MAC_5_641);
	MAC_5_642: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_642, data_out=>output_MAC_5_642);
	MAC_5_643: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_643, data_out=>output_MAC_5_643);
	MAC_5_644: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_644, data_out=>output_MAC_5_644);
	MAC_5_645: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_645, data_out=>output_MAC_5_645);
	MAC_5_646: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_646, data_out=>output_MAC_5_646);
	MAC_5_647: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_647, data_out=>output_MAC_5_647);
	MAC_5_648: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_648, data_out=>output_MAC_5_648);
	MAC_5_649: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_649, data_out=>output_MAC_5_649);
	MAC_5_650: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_650, data_out=>output_MAC_5_650);
	MAC_5_651: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_651, data_out=>output_MAC_5_651);
	MAC_5_652: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_652, data_out=>output_MAC_5_652);
	MAC_5_653: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_653, data_out=>output_MAC_5_653);
	MAC_5_654: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_654, data_out=>output_MAC_5_654);
	MAC_5_655: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_655, data_out=>output_MAC_5_655);
	MAC_5_656: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_656, data_out=>output_MAC_5_656);
	MAC_5_657: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_657, data_out=>output_MAC_5_657);
	MAC_5_658: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_658, data_out=>output_MAC_5_658);
	MAC_5_659: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_659, data_out=>output_MAC_5_659);
	MAC_5_660: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_660, data_out=>output_MAC_5_660);
	MAC_5_661: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_661, data_out=>output_MAC_5_661);
	MAC_5_662: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_662, data_out=>output_MAC_5_662);
	MAC_5_663: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_663, data_out=>output_MAC_5_663);
	MAC_5_664: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_664, data_out=>output_MAC_5_664);
	MAC_5_665: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_665, data_out=>output_MAC_5_665);
	MAC_5_666: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_666, data_out=>output_MAC_5_666);
	MAC_5_667: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_667, data_out=>output_MAC_5_667);
	MAC_5_668: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_668, data_out=>output_MAC_5_668);
	MAC_5_669: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_669, data_out=>output_MAC_5_669);
	MAC_5_670: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_670, data_out=>output_MAC_5_670);
	MAC_5_671: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_671, data_out=>output_MAC_5_671);
	MAC_5_672: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_672, data_out=>output_MAC_5_672);
	MAC_5_673: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_673, data_out=>output_MAC_5_673);
	MAC_5_674: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_674, data_out=>output_MAC_5_674);
	MAC_5_675: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_675, data_out=>output_MAC_5_675);
	MAC_5_676: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_676, data_out=>output_MAC_5_676);
	MAC_5_677: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_677, data_out=>output_MAC_5_677);
	MAC_5_678: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_678, data_out=>output_MAC_5_678);
	MAC_5_679: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_679, data_out=>output_MAC_5_679);
	MAC_5_680: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_680, data_out=>output_MAC_5_680);
	MAC_5_681: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_681, data_out=>output_MAC_5_681);
	MAC_5_682: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_682, data_out=>output_MAC_5_682);
	MAC_5_683: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_683, data_out=>output_MAC_5_683);
	MAC_5_684: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_684, data_out=>output_MAC_5_684);
	MAC_5_685: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_685, data_out=>output_MAC_5_685);
	MAC_5_686: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_686, data_out=>output_MAC_5_686);
	MAC_5_687: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_687, data_out=>output_MAC_5_687);
	MAC_5_688: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_688, data_out=>output_MAC_5_688);
	MAC_5_689: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_689, data_out=>output_MAC_5_689);
	MAC_5_690: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_690, data_out=>output_MAC_5_690);
	MAC_5_691: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_691, data_out=>output_MAC_5_691);
	MAC_5_692: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_692, data_out=>output_MAC_5_692);
	MAC_5_693: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_693, data_out=>output_MAC_5_693);
	MAC_5_694: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_694, data_out=>output_MAC_5_694);
	MAC_5_695: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_695, data_out=>output_MAC_5_695);
	MAC_5_696: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_696, data_out=>output_MAC_5_696);
	MAC_5_697: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_697, data_out=>output_MAC_5_697);
	MAC_5_698: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_698, data_out=>output_MAC_5_698);
	MAC_5_699: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_699, data_out=>output_MAC_5_699);
	MAC_5_700: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_700, data_out=>output_MAC_5_700);
	MAC_5_701: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_701, data_out=>output_MAC_5_701);
	MAC_5_702: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_702, data_out=>output_MAC_5_702);
	MAC_5_703: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_703, data_out=>output_MAC_5_703);
	MAC_5_704: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_704, data_out=>output_MAC_5_704);
	MAC_5_705: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_705, data_out=>output_MAC_5_705);
	MAC_5_706: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_706, data_out=>output_MAC_5_706);
	MAC_5_707: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_707, data_out=>output_MAC_5_707);
	MAC_5_708: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_708, data_out=>output_MAC_5_708);
	MAC_5_709: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_709, data_out=>output_MAC_5_709);
	MAC_5_710: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_710, data_out=>output_MAC_5_710);
	MAC_5_711: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_711, data_out=>output_MAC_5_711);
	MAC_5_712: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_712, data_out=>output_MAC_5_712);
	MAC_5_713: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_713, data_out=>output_MAC_5_713);
	MAC_5_714: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_714, data_out=>output_MAC_5_714);
	MAC_5_715: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_715, data_out=>output_MAC_5_715);
	MAC_5_716: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_716, data_out=>output_MAC_5_716);
	MAC_5_717: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_717, data_out=>output_MAC_5_717);
	MAC_5_718: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_718, data_out=>output_MAC_5_718);
	MAC_5_719: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_719, data_out=>output_MAC_5_719);
	MAC_5_720: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_720, data_out=>output_MAC_5_720);
	MAC_5_721: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_721, data_out=>output_MAC_5_721);
	MAC_5_722: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_722, data_out=>output_MAC_5_722);
	MAC_5_723: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_723, data_out=>output_MAC_5_723);
	MAC_5_724: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_724, data_out=>output_MAC_5_724);
	MAC_5_725: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_725, data_out=>output_MAC_5_725);
	MAC_5_726: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_726, data_out=>output_MAC_5_726);
	MAC_5_727: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_727, data_out=>output_MAC_5_727);
	MAC_5_728: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_728, data_out=>output_MAC_5_728);
	MAC_5_729: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_729, data_out=>output_MAC_5_729);
	MAC_5_730: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_730, data_out=>output_MAC_5_730);
	MAC_5_731: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_731, data_out=>output_MAC_5_731);
	MAC_5_732: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_732, data_out=>output_MAC_5_732);
	MAC_5_733: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_733, data_out=>output_MAC_5_733);
	MAC_5_734: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_734, data_out=>output_MAC_5_734);
	MAC_5_735: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_735, data_out=>output_MAC_5_735);
	MAC_5_736: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_736, data_out=>output_MAC_5_736);
	MAC_5_737: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_737, data_out=>output_MAC_5_737);
	MAC_5_738: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_738, data_out=>output_MAC_5_738);
	MAC_5_739: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_739, data_out=>output_MAC_5_739);
	MAC_5_740: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_740, data_out=>output_MAC_5_740);
	MAC_5_741: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_741, data_out=>output_MAC_5_741);
	MAC_5_742: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_742, data_out=>output_MAC_5_742);
	MAC_5_743: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_743, data_out=>output_MAC_5_743);
	MAC_5_744: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_744, data_out=>output_MAC_5_744);
	MAC_5_745: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_745, data_out=>output_MAC_5_745);
	MAC_5_746: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_746, data_out=>output_MAC_5_746);
	MAC_5_747: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_747, data_out=>output_MAC_5_747);
	MAC_5_748: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_748, data_out=>output_MAC_5_748);
	MAC_5_749: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_749, data_out=>output_MAC_5_749);
	MAC_5_750: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_750, data_out=>output_MAC_5_750);
	MAC_5_751: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_751, data_out=>output_MAC_5_751);
	MAC_5_752: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_752, data_out=>output_MAC_5_752);
	MAC_5_753: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_753, data_out=>output_MAC_5_753);
	MAC_5_754: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_754, data_out=>output_MAC_5_754);
	MAC_5_755: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_755, data_out=>output_MAC_5_755);
	MAC_5_756: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_756, data_out=>output_MAC_5_756);
	MAC_5_757: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_757, data_out=>output_MAC_5_757);
	MAC_5_758: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_758, data_out=>output_MAC_5_758);
	MAC_5_759: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_759, data_out=>output_MAC_5_759);
	MAC_5_760: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_760, data_out=>output_MAC_5_760);
	MAC_5_761: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_761, data_out=>output_MAC_5_761);
	MAC_5_762: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_762, data_out=>output_MAC_5_762);
	MAC_5_763: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_763, data_out=>output_MAC_5_763);
	MAC_5_764: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_764, data_out=>output_MAC_5_764);
	MAC_5_765: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_765, data_out=>output_MAC_5_765);
	MAC_5_766: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_766, data_out=>output_MAC_5_766);
	MAC_5_767: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_5, data_in_B=>input_col_767, data_out=>output_MAC_5_767);
	MAC_6_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_0, data_out=>output_MAC_6_0);
	MAC_6_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_1, data_out=>output_MAC_6_1);
	MAC_6_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_2, data_out=>output_MAC_6_2);
	MAC_6_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_3, data_out=>output_MAC_6_3);
	MAC_6_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_4, data_out=>output_MAC_6_4);
	MAC_6_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_5, data_out=>output_MAC_6_5);
	MAC_6_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_6, data_out=>output_MAC_6_6);
	MAC_6_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_7, data_out=>output_MAC_6_7);
	MAC_6_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_8, data_out=>output_MAC_6_8);
	MAC_6_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_9, data_out=>output_MAC_6_9);
	MAC_6_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_10, data_out=>output_MAC_6_10);
	MAC_6_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_11, data_out=>output_MAC_6_11);
	MAC_6_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_12, data_out=>output_MAC_6_12);
	MAC_6_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_13, data_out=>output_MAC_6_13);
	MAC_6_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_14, data_out=>output_MAC_6_14);
	MAC_6_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_15, data_out=>output_MAC_6_15);
	MAC_6_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_16, data_out=>output_MAC_6_16);
	MAC_6_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_17, data_out=>output_MAC_6_17);
	MAC_6_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_18, data_out=>output_MAC_6_18);
	MAC_6_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_19, data_out=>output_MAC_6_19);
	MAC_6_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_20, data_out=>output_MAC_6_20);
	MAC_6_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_21, data_out=>output_MAC_6_21);
	MAC_6_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_22, data_out=>output_MAC_6_22);
	MAC_6_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_23, data_out=>output_MAC_6_23);
	MAC_6_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_24, data_out=>output_MAC_6_24);
	MAC_6_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_25, data_out=>output_MAC_6_25);
	MAC_6_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_26, data_out=>output_MAC_6_26);
	MAC_6_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_27, data_out=>output_MAC_6_27);
	MAC_6_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_28, data_out=>output_MAC_6_28);
	MAC_6_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_29, data_out=>output_MAC_6_29);
	MAC_6_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_30, data_out=>output_MAC_6_30);
	MAC_6_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_31, data_out=>output_MAC_6_31);
	MAC_6_32: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_32, data_out=>output_MAC_6_32);
	MAC_6_33: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_33, data_out=>output_MAC_6_33);
	MAC_6_34: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_34, data_out=>output_MAC_6_34);
	MAC_6_35: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_35, data_out=>output_MAC_6_35);
	MAC_6_36: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_36, data_out=>output_MAC_6_36);
	MAC_6_37: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_37, data_out=>output_MAC_6_37);
	MAC_6_38: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_38, data_out=>output_MAC_6_38);
	MAC_6_39: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_39, data_out=>output_MAC_6_39);
	MAC_6_40: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_40, data_out=>output_MAC_6_40);
	MAC_6_41: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_41, data_out=>output_MAC_6_41);
	MAC_6_42: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_42, data_out=>output_MAC_6_42);
	MAC_6_43: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_43, data_out=>output_MAC_6_43);
	MAC_6_44: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_44, data_out=>output_MAC_6_44);
	MAC_6_45: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_45, data_out=>output_MAC_6_45);
	MAC_6_46: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_46, data_out=>output_MAC_6_46);
	MAC_6_47: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_47, data_out=>output_MAC_6_47);
	MAC_6_48: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_48, data_out=>output_MAC_6_48);
	MAC_6_49: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_49, data_out=>output_MAC_6_49);
	MAC_6_50: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_50, data_out=>output_MAC_6_50);
	MAC_6_51: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_51, data_out=>output_MAC_6_51);
	MAC_6_52: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_52, data_out=>output_MAC_6_52);
	MAC_6_53: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_53, data_out=>output_MAC_6_53);
	MAC_6_54: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_54, data_out=>output_MAC_6_54);
	MAC_6_55: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_55, data_out=>output_MAC_6_55);
	MAC_6_56: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_56, data_out=>output_MAC_6_56);
	MAC_6_57: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_57, data_out=>output_MAC_6_57);
	MAC_6_58: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_58, data_out=>output_MAC_6_58);
	MAC_6_59: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_59, data_out=>output_MAC_6_59);
	MAC_6_60: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_60, data_out=>output_MAC_6_60);
	MAC_6_61: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_61, data_out=>output_MAC_6_61);
	MAC_6_62: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_62, data_out=>output_MAC_6_62);
	MAC_6_63: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_63, data_out=>output_MAC_6_63);
	MAC_6_64: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_64, data_out=>output_MAC_6_64);
	MAC_6_65: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_65, data_out=>output_MAC_6_65);
	MAC_6_66: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_66, data_out=>output_MAC_6_66);
	MAC_6_67: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_67, data_out=>output_MAC_6_67);
	MAC_6_68: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_68, data_out=>output_MAC_6_68);
	MAC_6_69: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_69, data_out=>output_MAC_6_69);
	MAC_6_70: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_70, data_out=>output_MAC_6_70);
	MAC_6_71: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_71, data_out=>output_MAC_6_71);
	MAC_6_72: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_72, data_out=>output_MAC_6_72);
	MAC_6_73: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_73, data_out=>output_MAC_6_73);
	MAC_6_74: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_74, data_out=>output_MAC_6_74);
	MAC_6_75: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_75, data_out=>output_MAC_6_75);
	MAC_6_76: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_76, data_out=>output_MAC_6_76);
	MAC_6_77: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_77, data_out=>output_MAC_6_77);
	MAC_6_78: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_78, data_out=>output_MAC_6_78);
	MAC_6_79: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_79, data_out=>output_MAC_6_79);
	MAC_6_80: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_80, data_out=>output_MAC_6_80);
	MAC_6_81: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_81, data_out=>output_MAC_6_81);
	MAC_6_82: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_82, data_out=>output_MAC_6_82);
	MAC_6_83: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_83, data_out=>output_MAC_6_83);
	MAC_6_84: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_84, data_out=>output_MAC_6_84);
	MAC_6_85: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_85, data_out=>output_MAC_6_85);
	MAC_6_86: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_86, data_out=>output_MAC_6_86);
	MAC_6_87: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_87, data_out=>output_MAC_6_87);
	MAC_6_88: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_88, data_out=>output_MAC_6_88);
	MAC_6_89: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_89, data_out=>output_MAC_6_89);
	MAC_6_90: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_90, data_out=>output_MAC_6_90);
	MAC_6_91: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_91, data_out=>output_MAC_6_91);
	MAC_6_92: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_92, data_out=>output_MAC_6_92);
	MAC_6_93: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_93, data_out=>output_MAC_6_93);
	MAC_6_94: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_94, data_out=>output_MAC_6_94);
	MAC_6_95: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_95, data_out=>output_MAC_6_95);
	MAC_6_96: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_96, data_out=>output_MAC_6_96);
	MAC_6_97: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_97, data_out=>output_MAC_6_97);
	MAC_6_98: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_98, data_out=>output_MAC_6_98);
	MAC_6_99: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_99, data_out=>output_MAC_6_99);
	MAC_6_100: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_100, data_out=>output_MAC_6_100);
	MAC_6_101: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_101, data_out=>output_MAC_6_101);
	MAC_6_102: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_102, data_out=>output_MAC_6_102);
	MAC_6_103: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_103, data_out=>output_MAC_6_103);
	MAC_6_104: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_104, data_out=>output_MAC_6_104);
	MAC_6_105: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_105, data_out=>output_MAC_6_105);
	MAC_6_106: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_106, data_out=>output_MAC_6_106);
	MAC_6_107: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_107, data_out=>output_MAC_6_107);
	MAC_6_108: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_108, data_out=>output_MAC_6_108);
	MAC_6_109: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_109, data_out=>output_MAC_6_109);
	MAC_6_110: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_110, data_out=>output_MAC_6_110);
	MAC_6_111: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_111, data_out=>output_MAC_6_111);
	MAC_6_112: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_112, data_out=>output_MAC_6_112);
	MAC_6_113: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_113, data_out=>output_MAC_6_113);
	MAC_6_114: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_114, data_out=>output_MAC_6_114);
	MAC_6_115: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_115, data_out=>output_MAC_6_115);
	MAC_6_116: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_116, data_out=>output_MAC_6_116);
	MAC_6_117: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_117, data_out=>output_MAC_6_117);
	MAC_6_118: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_118, data_out=>output_MAC_6_118);
	MAC_6_119: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_119, data_out=>output_MAC_6_119);
	MAC_6_120: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_120, data_out=>output_MAC_6_120);
	MAC_6_121: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_121, data_out=>output_MAC_6_121);
	MAC_6_122: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_122, data_out=>output_MAC_6_122);
	MAC_6_123: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_123, data_out=>output_MAC_6_123);
	MAC_6_124: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_124, data_out=>output_MAC_6_124);
	MAC_6_125: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_125, data_out=>output_MAC_6_125);
	MAC_6_126: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_126, data_out=>output_MAC_6_126);
	MAC_6_127: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_127, data_out=>output_MAC_6_127);
	MAC_6_128: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_128, data_out=>output_MAC_6_128);
	MAC_6_129: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_129, data_out=>output_MAC_6_129);
	MAC_6_130: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_130, data_out=>output_MAC_6_130);
	MAC_6_131: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_131, data_out=>output_MAC_6_131);
	MAC_6_132: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_132, data_out=>output_MAC_6_132);
	MAC_6_133: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_133, data_out=>output_MAC_6_133);
	MAC_6_134: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_134, data_out=>output_MAC_6_134);
	MAC_6_135: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_135, data_out=>output_MAC_6_135);
	MAC_6_136: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_136, data_out=>output_MAC_6_136);
	MAC_6_137: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_137, data_out=>output_MAC_6_137);
	MAC_6_138: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_138, data_out=>output_MAC_6_138);
	MAC_6_139: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_139, data_out=>output_MAC_6_139);
	MAC_6_140: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_140, data_out=>output_MAC_6_140);
	MAC_6_141: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_141, data_out=>output_MAC_6_141);
	MAC_6_142: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_142, data_out=>output_MAC_6_142);
	MAC_6_143: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_143, data_out=>output_MAC_6_143);
	MAC_6_144: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_144, data_out=>output_MAC_6_144);
	MAC_6_145: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_145, data_out=>output_MAC_6_145);
	MAC_6_146: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_146, data_out=>output_MAC_6_146);
	MAC_6_147: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_147, data_out=>output_MAC_6_147);
	MAC_6_148: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_148, data_out=>output_MAC_6_148);
	MAC_6_149: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_149, data_out=>output_MAC_6_149);
	MAC_6_150: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_150, data_out=>output_MAC_6_150);
	MAC_6_151: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_151, data_out=>output_MAC_6_151);
	MAC_6_152: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_152, data_out=>output_MAC_6_152);
	MAC_6_153: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_153, data_out=>output_MAC_6_153);
	MAC_6_154: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_154, data_out=>output_MAC_6_154);
	MAC_6_155: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_155, data_out=>output_MAC_6_155);
	MAC_6_156: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_156, data_out=>output_MAC_6_156);
	MAC_6_157: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_157, data_out=>output_MAC_6_157);
	MAC_6_158: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_158, data_out=>output_MAC_6_158);
	MAC_6_159: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_159, data_out=>output_MAC_6_159);
	MAC_6_160: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_160, data_out=>output_MAC_6_160);
	MAC_6_161: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_161, data_out=>output_MAC_6_161);
	MAC_6_162: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_162, data_out=>output_MAC_6_162);
	MAC_6_163: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_163, data_out=>output_MAC_6_163);
	MAC_6_164: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_164, data_out=>output_MAC_6_164);
	MAC_6_165: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_165, data_out=>output_MAC_6_165);
	MAC_6_166: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_166, data_out=>output_MAC_6_166);
	MAC_6_167: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_167, data_out=>output_MAC_6_167);
	MAC_6_168: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_168, data_out=>output_MAC_6_168);
	MAC_6_169: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_169, data_out=>output_MAC_6_169);
	MAC_6_170: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_170, data_out=>output_MAC_6_170);
	MAC_6_171: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_171, data_out=>output_MAC_6_171);
	MAC_6_172: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_172, data_out=>output_MAC_6_172);
	MAC_6_173: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_173, data_out=>output_MAC_6_173);
	MAC_6_174: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_174, data_out=>output_MAC_6_174);
	MAC_6_175: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_175, data_out=>output_MAC_6_175);
	MAC_6_176: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_176, data_out=>output_MAC_6_176);
	MAC_6_177: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_177, data_out=>output_MAC_6_177);
	MAC_6_178: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_178, data_out=>output_MAC_6_178);
	MAC_6_179: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_179, data_out=>output_MAC_6_179);
	MAC_6_180: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_180, data_out=>output_MAC_6_180);
	MAC_6_181: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_181, data_out=>output_MAC_6_181);
	MAC_6_182: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_182, data_out=>output_MAC_6_182);
	MAC_6_183: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_183, data_out=>output_MAC_6_183);
	MAC_6_184: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_184, data_out=>output_MAC_6_184);
	MAC_6_185: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_185, data_out=>output_MAC_6_185);
	MAC_6_186: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_186, data_out=>output_MAC_6_186);
	MAC_6_187: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_187, data_out=>output_MAC_6_187);
	MAC_6_188: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_188, data_out=>output_MAC_6_188);
	MAC_6_189: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_189, data_out=>output_MAC_6_189);
	MAC_6_190: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_190, data_out=>output_MAC_6_190);
	MAC_6_191: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_191, data_out=>output_MAC_6_191);
	MAC_6_192: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_192, data_out=>output_MAC_6_192);
	MAC_6_193: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_193, data_out=>output_MAC_6_193);
	MAC_6_194: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_194, data_out=>output_MAC_6_194);
	MAC_6_195: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_195, data_out=>output_MAC_6_195);
	MAC_6_196: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_196, data_out=>output_MAC_6_196);
	MAC_6_197: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_197, data_out=>output_MAC_6_197);
	MAC_6_198: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_198, data_out=>output_MAC_6_198);
	MAC_6_199: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_199, data_out=>output_MAC_6_199);
	MAC_6_200: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_200, data_out=>output_MAC_6_200);
	MAC_6_201: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_201, data_out=>output_MAC_6_201);
	MAC_6_202: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_202, data_out=>output_MAC_6_202);
	MAC_6_203: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_203, data_out=>output_MAC_6_203);
	MAC_6_204: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_204, data_out=>output_MAC_6_204);
	MAC_6_205: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_205, data_out=>output_MAC_6_205);
	MAC_6_206: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_206, data_out=>output_MAC_6_206);
	MAC_6_207: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_207, data_out=>output_MAC_6_207);
	MAC_6_208: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_208, data_out=>output_MAC_6_208);
	MAC_6_209: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_209, data_out=>output_MAC_6_209);
	MAC_6_210: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_210, data_out=>output_MAC_6_210);
	MAC_6_211: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_211, data_out=>output_MAC_6_211);
	MAC_6_212: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_212, data_out=>output_MAC_6_212);
	MAC_6_213: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_213, data_out=>output_MAC_6_213);
	MAC_6_214: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_214, data_out=>output_MAC_6_214);
	MAC_6_215: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_215, data_out=>output_MAC_6_215);
	MAC_6_216: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_216, data_out=>output_MAC_6_216);
	MAC_6_217: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_217, data_out=>output_MAC_6_217);
	MAC_6_218: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_218, data_out=>output_MAC_6_218);
	MAC_6_219: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_219, data_out=>output_MAC_6_219);
	MAC_6_220: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_220, data_out=>output_MAC_6_220);
	MAC_6_221: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_221, data_out=>output_MAC_6_221);
	MAC_6_222: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_222, data_out=>output_MAC_6_222);
	MAC_6_223: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_223, data_out=>output_MAC_6_223);
	MAC_6_224: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_224, data_out=>output_MAC_6_224);
	MAC_6_225: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_225, data_out=>output_MAC_6_225);
	MAC_6_226: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_226, data_out=>output_MAC_6_226);
	MAC_6_227: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_227, data_out=>output_MAC_6_227);
	MAC_6_228: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_228, data_out=>output_MAC_6_228);
	MAC_6_229: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_229, data_out=>output_MAC_6_229);
	MAC_6_230: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_230, data_out=>output_MAC_6_230);
	MAC_6_231: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_231, data_out=>output_MAC_6_231);
	MAC_6_232: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_232, data_out=>output_MAC_6_232);
	MAC_6_233: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_233, data_out=>output_MAC_6_233);
	MAC_6_234: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_234, data_out=>output_MAC_6_234);
	MAC_6_235: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_235, data_out=>output_MAC_6_235);
	MAC_6_236: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_236, data_out=>output_MAC_6_236);
	MAC_6_237: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_237, data_out=>output_MAC_6_237);
	MAC_6_238: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_238, data_out=>output_MAC_6_238);
	MAC_6_239: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_239, data_out=>output_MAC_6_239);
	MAC_6_240: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_240, data_out=>output_MAC_6_240);
	MAC_6_241: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_241, data_out=>output_MAC_6_241);
	MAC_6_242: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_242, data_out=>output_MAC_6_242);
	MAC_6_243: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_243, data_out=>output_MAC_6_243);
	MAC_6_244: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_244, data_out=>output_MAC_6_244);
	MAC_6_245: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_245, data_out=>output_MAC_6_245);
	MAC_6_246: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_246, data_out=>output_MAC_6_246);
	MAC_6_247: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_247, data_out=>output_MAC_6_247);
	MAC_6_248: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_248, data_out=>output_MAC_6_248);
	MAC_6_249: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_249, data_out=>output_MAC_6_249);
	MAC_6_250: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_250, data_out=>output_MAC_6_250);
	MAC_6_251: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_251, data_out=>output_MAC_6_251);
	MAC_6_252: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_252, data_out=>output_MAC_6_252);
	MAC_6_253: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_253, data_out=>output_MAC_6_253);
	MAC_6_254: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_254, data_out=>output_MAC_6_254);
	MAC_6_255: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_255, data_out=>output_MAC_6_255);
	MAC_6_256: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_256, data_out=>output_MAC_6_256);
	MAC_6_257: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_257, data_out=>output_MAC_6_257);
	MAC_6_258: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_258, data_out=>output_MAC_6_258);
	MAC_6_259: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_259, data_out=>output_MAC_6_259);
	MAC_6_260: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_260, data_out=>output_MAC_6_260);
	MAC_6_261: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_261, data_out=>output_MAC_6_261);
	MAC_6_262: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_262, data_out=>output_MAC_6_262);
	MAC_6_263: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_263, data_out=>output_MAC_6_263);
	MAC_6_264: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_264, data_out=>output_MAC_6_264);
	MAC_6_265: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_265, data_out=>output_MAC_6_265);
	MAC_6_266: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_266, data_out=>output_MAC_6_266);
	MAC_6_267: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_267, data_out=>output_MAC_6_267);
	MAC_6_268: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_268, data_out=>output_MAC_6_268);
	MAC_6_269: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_269, data_out=>output_MAC_6_269);
	MAC_6_270: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_270, data_out=>output_MAC_6_270);
	MAC_6_271: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_271, data_out=>output_MAC_6_271);
	MAC_6_272: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_272, data_out=>output_MAC_6_272);
	MAC_6_273: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_273, data_out=>output_MAC_6_273);
	MAC_6_274: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_274, data_out=>output_MAC_6_274);
	MAC_6_275: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_275, data_out=>output_MAC_6_275);
	MAC_6_276: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_276, data_out=>output_MAC_6_276);
	MAC_6_277: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_277, data_out=>output_MAC_6_277);
	MAC_6_278: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_278, data_out=>output_MAC_6_278);
	MAC_6_279: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_279, data_out=>output_MAC_6_279);
	MAC_6_280: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_280, data_out=>output_MAC_6_280);
	MAC_6_281: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_281, data_out=>output_MAC_6_281);
	MAC_6_282: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_282, data_out=>output_MAC_6_282);
	MAC_6_283: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_283, data_out=>output_MAC_6_283);
	MAC_6_284: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_284, data_out=>output_MAC_6_284);
	MAC_6_285: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_285, data_out=>output_MAC_6_285);
	MAC_6_286: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_286, data_out=>output_MAC_6_286);
	MAC_6_287: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_287, data_out=>output_MAC_6_287);
	MAC_6_288: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_288, data_out=>output_MAC_6_288);
	MAC_6_289: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_289, data_out=>output_MAC_6_289);
	MAC_6_290: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_290, data_out=>output_MAC_6_290);
	MAC_6_291: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_291, data_out=>output_MAC_6_291);
	MAC_6_292: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_292, data_out=>output_MAC_6_292);
	MAC_6_293: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_293, data_out=>output_MAC_6_293);
	MAC_6_294: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_294, data_out=>output_MAC_6_294);
	MAC_6_295: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_295, data_out=>output_MAC_6_295);
	MAC_6_296: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_296, data_out=>output_MAC_6_296);
	MAC_6_297: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_297, data_out=>output_MAC_6_297);
	MAC_6_298: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_298, data_out=>output_MAC_6_298);
	MAC_6_299: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_299, data_out=>output_MAC_6_299);
	MAC_6_300: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_300, data_out=>output_MAC_6_300);
	MAC_6_301: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_301, data_out=>output_MAC_6_301);
	MAC_6_302: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_302, data_out=>output_MAC_6_302);
	MAC_6_303: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_303, data_out=>output_MAC_6_303);
	MAC_6_304: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_304, data_out=>output_MAC_6_304);
	MAC_6_305: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_305, data_out=>output_MAC_6_305);
	MAC_6_306: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_306, data_out=>output_MAC_6_306);
	MAC_6_307: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_307, data_out=>output_MAC_6_307);
	MAC_6_308: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_308, data_out=>output_MAC_6_308);
	MAC_6_309: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_309, data_out=>output_MAC_6_309);
	MAC_6_310: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_310, data_out=>output_MAC_6_310);
	MAC_6_311: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_311, data_out=>output_MAC_6_311);
	MAC_6_312: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_312, data_out=>output_MAC_6_312);
	MAC_6_313: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_313, data_out=>output_MAC_6_313);
	MAC_6_314: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_314, data_out=>output_MAC_6_314);
	MAC_6_315: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_315, data_out=>output_MAC_6_315);
	MAC_6_316: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_316, data_out=>output_MAC_6_316);
	MAC_6_317: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_317, data_out=>output_MAC_6_317);
	MAC_6_318: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_318, data_out=>output_MAC_6_318);
	MAC_6_319: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_319, data_out=>output_MAC_6_319);
	MAC_6_320: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_320, data_out=>output_MAC_6_320);
	MAC_6_321: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_321, data_out=>output_MAC_6_321);
	MAC_6_322: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_322, data_out=>output_MAC_6_322);
	MAC_6_323: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_323, data_out=>output_MAC_6_323);
	MAC_6_324: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_324, data_out=>output_MAC_6_324);
	MAC_6_325: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_325, data_out=>output_MAC_6_325);
	MAC_6_326: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_326, data_out=>output_MAC_6_326);
	MAC_6_327: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_327, data_out=>output_MAC_6_327);
	MAC_6_328: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_328, data_out=>output_MAC_6_328);
	MAC_6_329: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_329, data_out=>output_MAC_6_329);
	MAC_6_330: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_330, data_out=>output_MAC_6_330);
	MAC_6_331: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_331, data_out=>output_MAC_6_331);
	MAC_6_332: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_332, data_out=>output_MAC_6_332);
	MAC_6_333: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_333, data_out=>output_MAC_6_333);
	MAC_6_334: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_334, data_out=>output_MAC_6_334);
	MAC_6_335: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_335, data_out=>output_MAC_6_335);
	MAC_6_336: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_336, data_out=>output_MAC_6_336);
	MAC_6_337: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_337, data_out=>output_MAC_6_337);
	MAC_6_338: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_338, data_out=>output_MAC_6_338);
	MAC_6_339: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_339, data_out=>output_MAC_6_339);
	MAC_6_340: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_340, data_out=>output_MAC_6_340);
	MAC_6_341: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_341, data_out=>output_MAC_6_341);
	MAC_6_342: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_342, data_out=>output_MAC_6_342);
	MAC_6_343: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_343, data_out=>output_MAC_6_343);
	MAC_6_344: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_344, data_out=>output_MAC_6_344);
	MAC_6_345: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_345, data_out=>output_MAC_6_345);
	MAC_6_346: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_346, data_out=>output_MAC_6_346);
	MAC_6_347: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_347, data_out=>output_MAC_6_347);
	MAC_6_348: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_348, data_out=>output_MAC_6_348);
	MAC_6_349: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_349, data_out=>output_MAC_6_349);
	MAC_6_350: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_350, data_out=>output_MAC_6_350);
	MAC_6_351: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_351, data_out=>output_MAC_6_351);
	MAC_6_352: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_352, data_out=>output_MAC_6_352);
	MAC_6_353: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_353, data_out=>output_MAC_6_353);
	MAC_6_354: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_354, data_out=>output_MAC_6_354);
	MAC_6_355: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_355, data_out=>output_MAC_6_355);
	MAC_6_356: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_356, data_out=>output_MAC_6_356);
	MAC_6_357: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_357, data_out=>output_MAC_6_357);
	MAC_6_358: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_358, data_out=>output_MAC_6_358);
	MAC_6_359: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_359, data_out=>output_MAC_6_359);
	MAC_6_360: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_360, data_out=>output_MAC_6_360);
	MAC_6_361: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_361, data_out=>output_MAC_6_361);
	MAC_6_362: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_362, data_out=>output_MAC_6_362);
	MAC_6_363: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_363, data_out=>output_MAC_6_363);
	MAC_6_364: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_364, data_out=>output_MAC_6_364);
	MAC_6_365: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_365, data_out=>output_MAC_6_365);
	MAC_6_366: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_366, data_out=>output_MAC_6_366);
	MAC_6_367: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_367, data_out=>output_MAC_6_367);
	MAC_6_368: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_368, data_out=>output_MAC_6_368);
	MAC_6_369: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_369, data_out=>output_MAC_6_369);
	MAC_6_370: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_370, data_out=>output_MAC_6_370);
	MAC_6_371: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_371, data_out=>output_MAC_6_371);
	MAC_6_372: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_372, data_out=>output_MAC_6_372);
	MAC_6_373: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_373, data_out=>output_MAC_6_373);
	MAC_6_374: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_374, data_out=>output_MAC_6_374);
	MAC_6_375: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_375, data_out=>output_MAC_6_375);
	MAC_6_376: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_376, data_out=>output_MAC_6_376);
	MAC_6_377: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_377, data_out=>output_MAC_6_377);
	MAC_6_378: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_378, data_out=>output_MAC_6_378);
	MAC_6_379: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_379, data_out=>output_MAC_6_379);
	MAC_6_380: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_380, data_out=>output_MAC_6_380);
	MAC_6_381: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_381, data_out=>output_MAC_6_381);
	MAC_6_382: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_382, data_out=>output_MAC_6_382);
	MAC_6_383: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_383, data_out=>output_MAC_6_383);
	MAC_6_384: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_384, data_out=>output_MAC_6_384);
	MAC_6_385: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_385, data_out=>output_MAC_6_385);
	MAC_6_386: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_386, data_out=>output_MAC_6_386);
	MAC_6_387: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_387, data_out=>output_MAC_6_387);
	MAC_6_388: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_388, data_out=>output_MAC_6_388);
	MAC_6_389: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_389, data_out=>output_MAC_6_389);
	MAC_6_390: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_390, data_out=>output_MAC_6_390);
	MAC_6_391: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_391, data_out=>output_MAC_6_391);
	MAC_6_392: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_392, data_out=>output_MAC_6_392);
	MAC_6_393: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_393, data_out=>output_MAC_6_393);
	MAC_6_394: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_394, data_out=>output_MAC_6_394);
	MAC_6_395: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_395, data_out=>output_MAC_6_395);
	MAC_6_396: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_396, data_out=>output_MAC_6_396);
	MAC_6_397: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_397, data_out=>output_MAC_6_397);
	MAC_6_398: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_398, data_out=>output_MAC_6_398);
	MAC_6_399: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_399, data_out=>output_MAC_6_399);
	MAC_6_400: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_400, data_out=>output_MAC_6_400);
	MAC_6_401: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_401, data_out=>output_MAC_6_401);
	MAC_6_402: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_402, data_out=>output_MAC_6_402);
	MAC_6_403: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_403, data_out=>output_MAC_6_403);
	MAC_6_404: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_404, data_out=>output_MAC_6_404);
	MAC_6_405: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_405, data_out=>output_MAC_6_405);
	MAC_6_406: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_406, data_out=>output_MAC_6_406);
	MAC_6_407: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_407, data_out=>output_MAC_6_407);
	MAC_6_408: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_408, data_out=>output_MAC_6_408);
	MAC_6_409: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_409, data_out=>output_MAC_6_409);
	MAC_6_410: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_410, data_out=>output_MAC_6_410);
	MAC_6_411: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_411, data_out=>output_MAC_6_411);
	MAC_6_412: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_412, data_out=>output_MAC_6_412);
	MAC_6_413: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_413, data_out=>output_MAC_6_413);
	MAC_6_414: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_414, data_out=>output_MAC_6_414);
	MAC_6_415: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_415, data_out=>output_MAC_6_415);
	MAC_6_416: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_416, data_out=>output_MAC_6_416);
	MAC_6_417: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_417, data_out=>output_MAC_6_417);
	MAC_6_418: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_418, data_out=>output_MAC_6_418);
	MAC_6_419: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_419, data_out=>output_MAC_6_419);
	MAC_6_420: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_420, data_out=>output_MAC_6_420);
	MAC_6_421: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_421, data_out=>output_MAC_6_421);
	MAC_6_422: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_422, data_out=>output_MAC_6_422);
	MAC_6_423: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_423, data_out=>output_MAC_6_423);
	MAC_6_424: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_424, data_out=>output_MAC_6_424);
	MAC_6_425: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_425, data_out=>output_MAC_6_425);
	MAC_6_426: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_426, data_out=>output_MAC_6_426);
	MAC_6_427: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_427, data_out=>output_MAC_6_427);
	MAC_6_428: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_428, data_out=>output_MAC_6_428);
	MAC_6_429: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_429, data_out=>output_MAC_6_429);
	MAC_6_430: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_430, data_out=>output_MAC_6_430);
	MAC_6_431: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_431, data_out=>output_MAC_6_431);
	MAC_6_432: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_432, data_out=>output_MAC_6_432);
	MAC_6_433: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_433, data_out=>output_MAC_6_433);
	MAC_6_434: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_434, data_out=>output_MAC_6_434);
	MAC_6_435: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_435, data_out=>output_MAC_6_435);
	MAC_6_436: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_436, data_out=>output_MAC_6_436);
	MAC_6_437: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_437, data_out=>output_MAC_6_437);
	MAC_6_438: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_438, data_out=>output_MAC_6_438);
	MAC_6_439: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_439, data_out=>output_MAC_6_439);
	MAC_6_440: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_440, data_out=>output_MAC_6_440);
	MAC_6_441: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_441, data_out=>output_MAC_6_441);
	MAC_6_442: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_442, data_out=>output_MAC_6_442);
	MAC_6_443: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_443, data_out=>output_MAC_6_443);
	MAC_6_444: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_444, data_out=>output_MAC_6_444);
	MAC_6_445: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_445, data_out=>output_MAC_6_445);
	MAC_6_446: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_446, data_out=>output_MAC_6_446);
	MAC_6_447: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_447, data_out=>output_MAC_6_447);
	MAC_6_448: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_448, data_out=>output_MAC_6_448);
	MAC_6_449: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_449, data_out=>output_MAC_6_449);
	MAC_6_450: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_450, data_out=>output_MAC_6_450);
	MAC_6_451: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_451, data_out=>output_MAC_6_451);
	MAC_6_452: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_452, data_out=>output_MAC_6_452);
	MAC_6_453: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_453, data_out=>output_MAC_6_453);
	MAC_6_454: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_454, data_out=>output_MAC_6_454);
	MAC_6_455: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_455, data_out=>output_MAC_6_455);
	MAC_6_456: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_456, data_out=>output_MAC_6_456);
	MAC_6_457: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_457, data_out=>output_MAC_6_457);
	MAC_6_458: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_458, data_out=>output_MAC_6_458);
	MAC_6_459: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_459, data_out=>output_MAC_6_459);
	MAC_6_460: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_460, data_out=>output_MAC_6_460);
	MAC_6_461: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_461, data_out=>output_MAC_6_461);
	MAC_6_462: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_462, data_out=>output_MAC_6_462);
	MAC_6_463: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_463, data_out=>output_MAC_6_463);
	MAC_6_464: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_464, data_out=>output_MAC_6_464);
	MAC_6_465: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_465, data_out=>output_MAC_6_465);
	MAC_6_466: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_466, data_out=>output_MAC_6_466);
	MAC_6_467: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_467, data_out=>output_MAC_6_467);
	MAC_6_468: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_468, data_out=>output_MAC_6_468);
	MAC_6_469: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_469, data_out=>output_MAC_6_469);
	MAC_6_470: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_470, data_out=>output_MAC_6_470);
	MAC_6_471: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_471, data_out=>output_MAC_6_471);
	MAC_6_472: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_472, data_out=>output_MAC_6_472);
	MAC_6_473: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_473, data_out=>output_MAC_6_473);
	MAC_6_474: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_474, data_out=>output_MAC_6_474);
	MAC_6_475: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_475, data_out=>output_MAC_6_475);
	MAC_6_476: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_476, data_out=>output_MAC_6_476);
	MAC_6_477: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_477, data_out=>output_MAC_6_477);
	MAC_6_478: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_478, data_out=>output_MAC_6_478);
	MAC_6_479: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_479, data_out=>output_MAC_6_479);
	MAC_6_480: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_480, data_out=>output_MAC_6_480);
	MAC_6_481: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_481, data_out=>output_MAC_6_481);
	MAC_6_482: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_482, data_out=>output_MAC_6_482);
	MAC_6_483: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_483, data_out=>output_MAC_6_483);
	MAC_6_484: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_484, data_out=>output_MAC_6_484);
	MAC_6_485: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_485, data_out=>output_MAC_6_485);
	MAC_6_486: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_486, data_out=>output_MAC_6_486);
	MAC_6_487: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_487, data_out=>output_MAC_6_487);
	MAC_6_488: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_488, data_out=>output_MAC_6_488);
	MAC_6_489: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_489, data_out=>output_MAC_6_489);
	MAC_6_490: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_490, data_out=>output_MAC_6_490);
	MAC_6_491: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_491, data_out=>output_MAC_6_491);
	MAC_6_492: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_492, data_out=>output_MAC_6_492);
	MAC_6_493: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_493, data_out=>output_MAC_6_493);
	MAC_6_494: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_494, data_out=>output_MAC_6_494);
	MAC_6_495: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_495, data_out=>output_MAC_6_495);
	MAC_6_496: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_496, data_out=>output_MAC_6_496);
	MAC_6_497: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_497, data_out=>output_MAC_6_497);
	MAC_6_498: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_498, data_out=>output_MAC_6_498);
	MAC_6_499: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_499, data_out=>output_MAC_6_499);
	MAC_6_500: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_500, data_out=>output_MAC_6_500);
	MAC_6_501: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_501, data_out=>output_MAC_6_501);
	MAC_6_502: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_502, data_out=>output_MAC_6_502);
	MAC_6_503: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_503, data_out=>output_MAC_6_503);
	MAC_6_504: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_504, data_out=>output_MAC_6_504);
	MAC_6_505: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_505, data_out=>output_MAC_6_505);
	MAC_6_506: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_506, data_out=>output_MAC_6_506);
	MAC_6_507: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_507, data_out=>output_MAC_6_507);
	MAC_6_508: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_508, data_out=>output_MAC_6_508);
	MAC_6_509: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_509, data_out=>output_MAC_6_509);
	MAC_6_510: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_510, data_out=>output_MAC_6_510);
	MAC_6_511: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_511, data_out=>output_MAC_6_511);
	MAC_6_512: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_512, data_out=>output_MAC_6_512);
	MAC_6_513: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_513, data_out=>output_MAC_6_513);
	MAC_6_514: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_514, data_out=>output_MAC_6_514);
	MAC_6_515: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_515, data_out=>output_MAC_6_515);
	MAC_6_516: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_516, data_out=>output_MAC_6_516);
	MAC_6_517: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_517, data_out=>output_MAC_6_517);
	MAC_6_518: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_518, data_out=>output_MAC_6_518);
	MAC_6_519: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_519, data_out=>output_MAC_6_519);
	MAC_6_520: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_520, data_out=>output_MAC_6_520);
	MAC_6_521: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_521, data_out=>output_MAC_6_521);
	MAC_6_522: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_522, data_out=>output_MAC_6_522);
	MAC_6_523: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_523, data_out=>output_MAC_6_523);
	MAC_6_524: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_524, data_out=>output_MAC_6_524);
	MAC_6_525: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_525, data_out=>output_MAC_6_525);
	MAC_6_526: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_526, data_out=>output_MAC_6_526);
	MAC_6_527: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_527, data_out=>output_MAC_6_527);
	MAC_6_528: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_528, data_out=>output_MAC_6_528);
	MAC_6_529: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_529, data_out=>output_MAC_6_529);
	MAC_6_530: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_530, data_out=>output_MAC_6_530);
	MAC_6_531: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_531, data_out=>output_MAC_6_531);
	MAC_6_532: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_532, data_out=>output_MAC_6_532);
	MAC_6_533: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_533, data_out=>output_MAC_6_533);
	MAC_6_534: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_534, data_out=>output_MAC_6_534);
	MAC_6_535: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_535, data_out=>output_MAC_6_535);
	MAC_6_536: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_536, data_out=>output_MAC_6_536);
	MAC_6_537: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_537, data_out=>output_MAC_6_537);
	MAC_6_538: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_538, data_out=>output_MAC_6_538);
	MAC_6_539: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_539, data_out=>output_MAC_6_539);
	MAC_6_540: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_540, data_out=>output_MAC_6_540);
	MAC_6_541: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_541, data_out=>output_MAC_6_541);
	MAC_6_542: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_542, data_out=>output_MAC_6_542);
	MAC_6_543: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_543, data_out=>output_MAC_6_543);
	MAC_6_544: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_544, data_out=>output_MAC_6_544);
	MAC_6_545: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_545, data_out=>output_MAC_6_545);
	MAC_6_546: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_546, data_out=>output_MAC_6_546);
	MAC_6_547: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_547, data_out=>output_MAC_6_547);
	MAC_6_548: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_548, data_out=>output_MAC_6_548);
	MAC_6_549: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_549, data_out=>output_MAC_6_549);
	MAC_6_550: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_550, data_out=>output_MAC_6_550);
	MAC_6_551: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_551, data_out=>output_MAC_6_551);
	MAC_6_552: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_552, data_out=>output_MAC_6_552);
	MAC_6_553: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_553, data_out=>output_MAC_6_553);
	MAC_6_554: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_554, data_out=>output_MAC_6_554);
	MAC_6_555: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_555, data_out=>output_MAC_6_555);
	MAC_6_556: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_556, data_out=>output_MAC_6_556);
	MAC_6_557: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_557, data_out=>output_MAC_6_557);
	MAC_6_558: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_558, data_out=>output_MAC_6_558);
	MAC_6_559: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_559, data_out=>output_MAC_6_559);
	MAC_6_560: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_560, data_out=>output_MAC_6_560);
	MAC_6_561: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_561, data_out=>output_MAC_6_561);
	MAC_6_562: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_562, data_out=>output_MAC_6_562);
	MAC_6_563: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_563, data_out=>output_MAC_6_563);
	MAC_6_564: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_564, data_out=>output_MAC_6_564);
	MAC_6_565: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_565, data_out=>output_MAC_6_565);
	MAC_6_566: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_566, data_out=>output_MAC_6_566);
	MAC_6_567: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_567, data_out=>output_MAC_6_567);
	MAC_6_568: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_568, data_out=>output_MAC_6_568);
	MAC_6_569: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_569, data_out=>output_MAC_6_569);
	MAC_6_570: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_570, data_out=>output_MAC_6_570);
	MAC_6_571: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_571, data_out=>output_MAC_6_571);
	MAC_6_572: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_572, data_out=>output_MAC_6_572);
	MAC_6_573: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_573, data_out=>output_MAC_6_573);
	MAC_6_574: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_574, data_out=>output_MAC_6_574);
	MAC_6_575: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_575, data_out=>output_MAC_6_575);
	MAC_6_576: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_576, data_out=>output_MAC_6_576);
	MAC_6_577: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_577, data_out=>output_MAC_6_577);
	MAC_6_578: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_578, data_out=>output_MAC_6_578);
	MAC_6_579: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_579, data_out=>output_MAC_6_579);
	MAC_6_580: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_580, data_out=>output_MAC_6_580);
	MAC_6_581: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_581, data_out=>output_MAC_6_581);
	MAC_6_582: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_582, data_out=>output_MAC_6_582);
	MAC_6_583: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_583, data_out=>output_MAC_6_583);
	MAC_6_584: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_584, data_out=>output_MAC_6_584);
	MAC_6_585: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_585, data_out=>output_MAC_6_585);
	MAC_6_586: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_586, data_out=>output_MAC_6_586);
	MAC_6_587: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_587, data_out=>output_MAC_6_587);
	MAC_6_588: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_588, data_out=>output_MAC_6_588);
	MAC_6_589: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_589, data_out=>output_MAC_6_589);
	MAC_6_590: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_590, data_out=>output_MAC_6_590);
	MAC_6_591: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_591, data_out=>output_MAC_6_591);
	MAC_6_592: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_592, data_out=>output_MAC_6_592);
	MAC_6_593: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_593, data_out=>output_MAC_6_593);
	MAC_6_594: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_594, data_out=>output_MAC_6_594);
	MAC_6_595: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_595, data_out=>output_MAC_6_595);
	MAC_6_596: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_596, data_out=>output_MAC_6_596);
	MAC_6_597: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_597, data_out=>output_MAC_6_597);
	MAC_6_598: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_598, data_out=>output_MAC_6_598);
	MAC_6_599: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_599, data_out=>output_MAC_6_599);
	MAC_6_600: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_600, data_out=>output_MAC_6_600);
	MAC_6_601: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_601, data_out=>output_MAC_6_601);
	MAC_6_602: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_602, data_out=>output_MAC_6_602);
	MAC_6_603: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_603, data_out=>output_MAC_6_603);
	MAC_6_604: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_604, data_out=>output_MAC_6_604);
	MAC_6_605: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_605, data_out=>output_MAC_6_605);
	MAC_6_606: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_606, data_out=>output_MAC_6_606);
	MAC_6_607: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_607, data_out=>output_MAC_6_607);
	MAC_6_608: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_608, data_out=>output_MAC_6_608);
	MAC_6_609: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_609, data_out=>output_MAC_6_609);
	MAC_6_610: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_610, data_out=>output_MAC_6_610);
	MAC_6_611: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_611, data_out=>output_MAC_6_611);
	MAC_6_612: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_612, data_out=>output_MAC_6_612);
	MAC_6_613: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_613, data_out=>output_MAC_6_613);
	MAC_6_614: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_614, data_out=>output_MAC_6_614);
	MAC_6_615: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_615, data_out=>output_MAC_6_615);
	MAC_6_616: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_616, data_out=>output_MAC_6_616);
	MAC_6_617: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_617, data_out=>output_MAC_6_617);
	MAC_6_618: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_618, data_out=>output_MAC_6_618);
	MAC_6_619: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_619, data_out=>output_MAC_6_619);
	MAC_6_620: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_620, data_out=>output_MAC_6_620);
	MAC_6_621: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_621, data_out=>output_MAC_6_621);
	MAC_6_622: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_622, data_out=>output_MAC_6_622);
	MAC_6_623: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_623, data_out=>output_MAC_6_623);
	MAC_6_624: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_624, data_out=>output_MAC_6_624);
	MAC_6_625: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_625, data_out=>output_MAC_6_625);
	MAC_6_626: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_626, data_out=>output_MAC_6_626);
	MAC_6_627: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_627, data_out=>output_MAC_6_627);
	MAC_6_628: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_628, data_out=>output_MAC_6_628);
	MAC_6_629: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_629, data_out=>output_MAC_6_629);
	MAC_6_630: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_630, data_out=>output_MAC_6_630);
	MAC_6_631: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_631, data_out=>output_MAC_6_631);
	MAC_6_632: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_632, data_out=>output_MAC_6_632);
	MAC_6_633: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_633, data_out=>output_MAC_6_633);
	MAC_6_634: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_634, data_out=>output_MAC_6_634);
	MAC_6_635: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_635, data_out=>output_MAC_6_635);
	MAC_6_636: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_636, data_out=>output_MAC_6_636);
	MAC_6_637: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_637, data_out=>output_MAC_6_637);
	MAC_6_638: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_638, data_out=>output_MAC_6_638);
	MAC_6_639: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_639, data_out=>output_MAC_6_639);
	MAC_6_640: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_640, data_out=>output_MAC_6_640);
	MAC_6_641: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_641, data_out=>output_MAC_6_641);
	MAC_6_642: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_642, data_out=>output_MAC_6_642);
	MAC_6_643: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_643, data_out=>output_MAC_6_643);
	MAC_6_644: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_644, data_out=>output_MAC_6_644);
	MAC_6_645: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_645, data_out=>output_MAC_6_645);
	MAC_6_646: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_646, data_out=>output_MAC_6_646);
	MAC_6_647: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_647, data_out=>output_MAC_6_647);
	MAC_6_648: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_648, data_out=>output_MAC_6_648);
	MAC_6_649: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_649, data_out=>output_MAC_6_649);
	MAC_6_650: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_650, data_out=>output_MAC_6_650);
	MAC_6_651: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_651, data_out=>output_MAC_6_651);
	MAC_6_652: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_652, data_out=>output_MAC_6_652);
	MAC_6_653: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_653, data_out=>output_MAC_6_653);
	MAC_6_654: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_654, data_out=>output_MAC_6_654);
	MAC_6_655: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_655, data_out=>output_MAC_6_655);
	MAC_6_656: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_656, data_out=>output_MAC_6_656);
	MAC_6_657: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_657, data_out=>output_MAC_6_657);
	MAC_6_658: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_658, data_out=>output_MAC_6_658);
	MAC_6_659: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_659, data_out=>output_MAC_6_659);
	MAC_6_660: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_660, data_out=>output_MAC_6_660);
	MAC_6_661: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_661, data_out=>output_MAC_6_661);
	MAC_6_662: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_662, data_out=>output_MAC_6_662);
	MAC_6_663: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_663, data_out=>output_MAC_6_663);
	MAC_6_664: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_664, data_out=>output_MAC_6_664);
	MAC_6_665: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_665, data_out=>output_MAC_6_665);
	MAC_6_666: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_666, data_out=>output_MAC_6_666);
	MAC_6_667: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_667, data_out=>output_MAC_6_667);
	MAC_6_668: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_668, data_out=>output_MAC_6_668);
	MAC_6_669: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_669, data_out=>output_MAC_6_669);
	MAC_6_670: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_670, data_out=>output_MAC_6_670);
	MAC_6_671: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_671, data_out=>output_MAC_6_671);
	MAC_6_672: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_672, data_out=>output_MAC_6_672);
	MAC_6_673: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_673, data_out=>output_MAC_6_673);
	MAC_6_674: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_674, data_out=>output_MAC_6_674);
	MAC_6_675: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_675, data_out=>output_MAC_6_675);
	MAC_6_676: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_676, data_out=>output_MAC_6_676);
	MAC_6_677: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_677, data_out=>output_MAC_6_677);
	MAC_6_678: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_678, data_out=>output_MAC_6_678);
	MAC_6_679: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_679, data_out=>output_MAC_6_679);
	MAC_6_680: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_680, data_out=>output_MAC_6_680);
	MAC_6_681: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_681, data_out=>output_MAC_6_681);
	MAC_6_682: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_682, data_out=>output_MAC_6_682);
	MAC_6_683: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_683, data_out=>output_MAC_6_683);
	MAC_6_684: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_684, data_out=>output_MAC_6_684);
	MAC_6_685: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_685, data_out=>output_MAC_6_685);
	MAC_6_686: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_686, data_out=>output_MAC_6_686);
	MAC_6_687: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_687, data_out=>output_MAC_6_687);
	MAC_6_688: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_688, data_out=>output_MAC_6_688);
	MAC_6_689: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_689, data_out=>output_MAC_6_689);
	MAC_6_690: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_690, data_out=>output_MAC_6_690);
	MAC_6_691: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_691, data_out=>output_MAC_6_691);
	MAC_6_692: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_692, data_out=>output_MAC_6_692);
	MAC_6_693: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_693, data_out=>output_MAC_6_693);
	MAC_6_694: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_694, data_out=>output_MAC_6_694);
	MAC_6_695: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_695, data_out=>output_MAC_6_695);
	MAC_6_696: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_696, data_out=>output_MAC_6_696);
	MAC_6_697: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_697, data_out=>output_MAC_6_697);
	MAC_6_698: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_698, data_out=>output_MAC_6_698);
	MAC_6_699: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_699, data_out=>output_MAC_6_699);
	MAC_6_700: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_700, data_out=>output_MAC_6_700);
	MAC_6_701: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_701, data_out=>output_MAC_6_701);
	MAC_6_702: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_702, data_out=>output_MAC_6_702);
	MAC_6_703: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_703, data_out=>output_MAC_6_703);
	MAC_6_704: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_704, data_out=>output_MAC_6_704);
	MAC_6_705: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_705, data_out=>output_MAC_6_705);
	MAC_6_706: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_706, data_out=>output_MAC_6_706);
	MAC_6_707: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_707, data_out=>output_MAC_6_707);
	MAC_6_708: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_708, data_out=>output_MAC_6_708);
	MAC_6_709: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_709, data_out=>output_MAC_6_709);
	MAC_6_710: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_710, data_out=>output_MAC_6_710);
	MAC_6_711: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_711, data_out=>output_MAC_6_711);
	MAC_6_712: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_712, data_out=>output_MAC_6_712);
	MAC_6_713: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_713, data_out=>output_MAC_6_713);
	MAC_6_714: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_714, data_out=>output_MAC_6_714);
	MAC_6_715: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_715, data_out=>output_MAC_6_715);
	MAC_6_716: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_716, data_out=>output_MAC_6_716);
	MAC_6_717: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_717, data_out=>output_MAC_6_717);
	MAC_6_718: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_718, data_out=>output_MAC_6_718);
	MAC_6_719: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_719, data_out=>output_MAC_6_719);
	MAC_6_720: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_720, data_out=>output_MAC_6_720);
	MAC_6_721: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_721, data_out=>output_MAC_6_721);
	MAC_6_722: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_722, data_out=>output_MAC_6_722);
	MAC_6_723: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_723, data_out=>output_MAC_6_723);
	MAC_6_724: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_724, data_out=>output_MAC_6_724);
	MAC_6_725: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_725, data_out=>output_MAC_6_725);
	MAC_6_726: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_726, data_out=>output_MAC_6_726);
	MAC_6_727: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_727, data_out=>output_MAC_6_727);
	MAC_6_728: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_728, data_out=>output_MAC_6_728);
	MAC_6_729: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_729, data_out=>output_MAC_6_729);
	MAC_6_730: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_730, data_out=>output_MAC_6_730);
	MAC_6_731: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_731, data_out=>output_MAC_6_731);
	MAC_6_732: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_732, data_out=>output_MAC_6_732);
	MAC_6_733: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_733, data_out=>output_MAC_6_733);
	MAC_6_734: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_734, data_out=>output_MAC_6_734);
	MAC_6_735: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_735, data_out=>output_MAC_6_735);
	MAC_6_736: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_736, data_out=>output_MAC_6_736);
	MAC_6_737: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_737, data_out=>output_MAC_6_737);
	MAC_6_738: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_738, data_out=>output_MAC_6_738);
	MAC_6_739: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_739, data_out=>output_MAC_6_739);
	MAC_6_740: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_740, data_out=>output_MAC_6_740);
	MAC_6_741: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_741, data_out=>output_MAC_6_741);
	MAC_6_742: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_742, data_out=>output_MAC_6_742);
	MAC_6_743: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_743, data_out=>output_MAC_6_743);
	MAC_6_744: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_744, data_out=>output_MAC_6_744);
	MAC_6_745: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_745, data_out=>output_MAC_6_745);
	MAC_6_746: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_746, data_out=>output_MAC_6_746);
	MAC_6_747: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_747, data_out=>output_MAC_6_747);
	MAC_6_748: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_748, data_out=>output_MAC_6_748);
	MAC_6_749: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_749, data_out=>output_MAC_6_749);
	MAC_6_750: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_750, data_out=>output_MAC_6_750);
	MAC_6_751: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_751, data_out=>output_MAC_6_751);
	MAC_6_752: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_752, data_out=>output_MAC_6_752);
	MAC_6_753: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_753, data_out=>output_MAC_6_753);
	MAC_6_754: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_754, data_out=>output_MAC_6_754);
	MAC_6_755: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_755, data_out=>output_MAC_6_755);
	MAC_6_756: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_756, data_out=>output_MAC_6_756);
	MAC_6_757: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_757, data_out=>output_MAC_6_757);
	MAC_6_758: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_758, data_out=>output_MAC_6_758);
	MAC_6_759: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_759, data_out=>output_MAC_6_759);
	MAC_6_760: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_760, data_out=>output_MAC_6_760);
	MAC_6_761: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_761, data_out=>output_MAC_6_761);
	MAC_6_762: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_762, data_out=>output_MAC_6_762);
	MAC_6_763: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_763, data_out=>output_MAC_6_763);
	MAC_6_764: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_764, data_out=>output_MAC_6_764);
	MAC_6_765: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_765, data_out=>output_MAC_6_765);
	MAC_6_766: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_766, data_out=>output_MAC_6_766);
	MAC_6_767: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_6, data_in_B=>input_col_767, data_out=>output_MAC_6_767);
	MAC_7_0: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_0, data_out=>output_MAC_7_0);
	MAC_7_1: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_1, data_out=>output_MAC_7_1);
	MAC_7_2: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_2, data_out=>output_MAC_7_2);
	MAC_7_3: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_3, data_out=>output_MAC_7_3);
	MAC_7_4: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_4, data_out=>output_MAC_7_4);
	MAC_7_5: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_5, data_out=>output_MAC_7_5);
	MAC_7_6: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_6, data_out=>output_MAC_7_6);
	MAC_7_7: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_7, data_out=>output_MAC_7_7);
	MAC_7_8: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_8, data_out=>output_MAC_7_8);
	MAC_7_9: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_9, data_out=>output_MAC_7_9);
	MAC_7_10: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_10, data_out=>output_MAC_7_10);
	MAC_7_11: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_11, data_out=>output_MAC_7_11);
	MAC_7_12: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_12, data_out=>output_MAC_7_12);
	MAC_7_13: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_13, data_out=>output_MAC_7_13);
	MAC_7_14: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_14, data_out=>output_MAC_7_14);
	MAC_7_15: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_15, data_out=>output_MAC_7_15);
	MAC_7_16: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_16, data_out=>output_MAC_7_16);
	MAC_7_17: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_17, data_out=>output_MAC_7_17);
	MAC_7_18: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_18, data_out=>output_MAC_7_18);
	MAC_7_19: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_19, data_out=>output_MAC_7_19);
	MAC_7_20: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_20, data_out=>output_MAC_7_20);
	MAC_7_21: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_21, data_out=>output_MAC_7_21);
	MAC_7_22: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_22, data_out=>output_MAC_7_22);
	MAC_7_23: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_23, data_out=>output_MAC_7_23);
	MAC_7_24: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_24, data_out=>output_MAC_7_24);
	MAC_7_25: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_25, data_out=>output_MAC_7_25);
	MAC_7_26: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_26, data_out=>output_MAC_7_26);
	MAC_7_27: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_27, data_out=>output_MAC_7_27);
	MAC_7_28: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_28, data_out=>output_MAC_7_28);
	MAC_7_29: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_29, data_out=>output_MAC_7_29);
	MAC_7_30: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_30, data_out=>output_MAC_7_30);
	MAC_7_31: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_31, data_out=>output_MAC_7_31);
	MAC_7_32: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_32, data_out=>output_MAC_7_32);
	MAC_7_33: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_33, data_out=>output_MAC_7_33);
	MAC_7_34: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_34, data_out=>output_MAC_7_34);
	MAC_7_35: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_35, data_out=>output_MAC_7_35);
	MAC_7_36: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_36, data_out=>output_MAC_7_36);
	MAC_7_37: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_37, data_out=>output_MAC_7_37);
	MAC_7_38: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_38, data_out=>output_MAC_7_38);
	MAC_7_39: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_39, data_out=>output_MAC_7_39);
	MAC_7_40: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_40, data_out=>output_MAC_7_40);
	MAC_7_41: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_41, data_out=>output_MAC_7_41);
	MAC_7_42: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_42, data_out=>output_MAC_7_42);
	MAC_7_43: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_43, data_out=>output_MAC_7_43);
	MAC_7_44: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_44, data_out=>output_MAC_7_44);
	MAC_7_45: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_45, data_out=>output_MAC_7_45);
	MAC_7_46: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_46, data_out=>output_MAC_7_46);
	MAC_7_47: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_47, data_out=>output_MAC_7_47);
	MAC_7_48: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_48, data_out=>output_MAC_7_48);
	MAC_7_49: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_49, data_out=>output_MAC_7_49);
	MAC_7_50: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_50, data_out=>output_MAC_7_50);
	MAC_7_51: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_51, data_out=>output_MAC_7_51);
	MAC_7_52: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_52, data_out=>output_MAC_7_52);
	MAC_7_53: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_53, data_out=>output_MAC_7_53);
	MAC_7_54: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_54, data_out=>output_MAC_7_54);
	MAC_7_55: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_55, data_out=>output_MAC_7_55);
	MAC_7_56: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_56, data_out=>output_MAC_7_56);
	MAC_7_57: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_57, data_out=>output_MAC_7_57);
	MAC_7_58: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_58, data_out=>output_MAC_7_58);
	MAC_7_59: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_59, data_out=>output_MAC_7_59);
	MAC_7_60: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_60, data_out=>output_MAC_7_60);
	MAC_7_61: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_61, data_out=>output_MAC_7_61);
	MAC_7_62: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_62, data_out=>output_MAC_7_62);
	MAC_7_63: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_63, data_out=>output_MAC_7_63);
	MAC_7_64: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_64, data_out=>output_MAC_7_64);
	MAC_7_65: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_65, data_out=>output_MAC_7_65);
	MAC_7_66: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_66, data_out=>output_MAC_7_66);
	MAC_7_67: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_67, data_out=>output_MAC_7_67);
	MAC_7_68: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_68, data_out=>output_MAC_7_68);
	MAC_7_69: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_69, data_out=>output_MAC_7_69);
	MAC_7_70: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_70, data_out=>output_MAC_7_70);
	MAC_7_71: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_71, data_out=>output_MAC_7_71);
	MAC_7_72: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_72, data_out=>output_MAC_7_72);
	MAC_7_73: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_73, data_out=>output_MAC_7_73);
	MAC_7_74: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_74, data_out=>output_MAC_7_74);
	MAC_7_75: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_75, data_out=>output_MAC_7_75);
	MAC_7_76: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_76, data_out=>output_MAC_7_76);
	MAC_7_77: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_77, data_out=>output_MAC_7_77);
	MAC_7_78: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_78, data_out=>output_MAC_7_78);
	MAC_7_79: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_79, data_out=>output_MAC_7_79);
	MAC_7_80: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_80, data_out=>output_MAC_7_80);
	MAC_7_81: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_81, data_out=>output_MAC_7_81);
	MAC_7_82: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_82, data_out=>output_MAC_7_82);
	MAC_7_83: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_83, data_out=>output_MAC_7_83);
	MAC_7_84: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_84, data_out=>output_MAC_7_84);
	MAC_7_85: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_85, data_out=>output_MAC_7_85);
	MAC_7_86: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_86, data_out=>output_MAC_7_86);
	MAC_7_87: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_87, data_out=>output_MAC_7_87);
	MAC_7_88: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_88, data_out=>output_MAC_7_88);
	MAC_7_89: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_89, data_out=>output_MAC_7_89);
	MAC_7_90: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_90, data_out=>output_MAC_7_90);
	MAC_7_91: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_91, data_out=>output_MAC_7_91);
	MAC_7_92: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_92, data_out=>output_MAC_7_92);
	MAC_7_93: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_93, data_out=>output_MAC_7_93);
	MAC_7_94: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_94, data_out=>output_MAC_7_94);
	MAC_7_95: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_95, data_out=>output_MAC_7_95);
	MAC_7_96: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_96, data_out=>output_MAC_7_96);
	MAC_7_97: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_97, data_out=>output_MAC_7_97);
	MAC_7_98: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_98, data_out=>output_MAC_7_98);
	MAC_7_99: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_99, data_out=>output_MAC_7_99);
	MAC_7_100: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_100, data_out=>output_MAC_7_100);
	MAC_7_101: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_101, data_out=>output_MAC_7_101);
	MAC_7_102: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_102, data_out=>output_MAC_7_102);
	MAC_7_103: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_103, data_out=>output_MAC_7_103);
	MAC_7_104: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_104, data_out=>output_MAC_7_104);
	MAC_7_105: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_105, data_out=>output_MAC_7_105);
	MAC_7_106: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_106, data_out=>output_MAC_7_106);
	MAC_7_107: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_107, data_out=>output_MAC_7_107);
	MAC_7_108: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_108, data_out=>output_MAC_7_108);
	MAC_7_109: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_109, data_out=>output_MAC_7_109);
	MAC_7_110: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_110, data_out=>output_MAC_7_110);
	MAC_7_111: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_111, data_out=>output_MAC_7_111);
	MAC_7_112: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_112, data_out=>output_MAC_7_112);
	MAC_7_113: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_113, data_out=>output_MAC_7_113);
	MAC_7_114: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_114, data_out=>output_MAC_7_114);
	MAC_7_115: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_115, data_out=>output_MAC_7_115);
	MAC_7_116: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_116, data_out=>output_MAC_7_116);
	MAC_7_117: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_117, data_out=>output_MAC_7_117);
	MAC_7_118: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_118, data_out=>output_MAC_7_118);
	MAC_7_119: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_119, data_out=>output_MAC_7_119);
	MAC_7_120: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_120, data_out=>output_MAC_7_120);
	MAC_7_121: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_121, data_out=>output_MAC_7_121);
	MAC_7_122: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_122, data_out=>output_MAC_7_122);
	MAC_7_123: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_123, data_out=>output_MAC_7_123);
	MAC_7_124: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_124, data_out=>output_MAC_7_124);
	MAC_7_125: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_125, data_out=>output_MAC_7_125);
	MAC_7_126: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_126, data_out=>output_MAC_7_126);
	MAC_7_127: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_127, data_out=>output_MAC_7_127);
	MAC_7_128: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_128, data_out=>output_MAC_7_128);
	MAC_7_129: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_129, data_out=>output_MAC_7_129);
	MAC_7_130: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_130, data_out=>output_MAC_7_130);
	MAC_7_131: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_131, data_out=>output_MAC_7_131);
	MAC_7_132: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_132, data_out=>output_MAC_7_132);
	MAC_7_133: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_133, data_out=>output_MAC_7_133);
	MAC_7_134: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_134, data_out=>output_MAC_7_134);
	MAC_7_135: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_135, data_out=>output_MAC_7_135);
	MAC_7_136: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_136, data_out=>output_MAC_7_136);
	MAC_7_137: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_137, data_out=>output_MAC_7_137);
	MAC_7_138: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_138, data_out=>output_MAC_7_138);
	MAC_7_139: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_139, data_out=>output_MAC_7_139);
	MAC_7_140: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_140, data_out=>output_MAC_7_140);
	MAC_7_141: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_141, data_out=>output_MAC_7_141);
	MAC_7_142: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_142, data_out=>output_MAC_7_142);
	MAC_7_143: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_143, data_out=>output_MAC_7_143);
	MAC_7_144: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_144, data_out=>output_MAC_7_144);
	MAC_7_145: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_145, data_out=>output_MAC_7_145);
	MAC_7_146: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_146, data_out=>output_MAC_7_146);
	MAC_7_147: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_147, data_out=>output_MAC_7_147);
	MAC_7_148: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_148, data_out=>output_MAC_7_148);
	MAC_7_149: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_149, data_out=>output_MAC_7_149);
	MAC_7_150: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_150, data_out=>output_MAC_7_150);
	MAC_7_151: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_151, data_out=>output_MAC_7_151);
	MAC_7_152: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_152, data_out=>output_MAC_7_152);
	MAC_7_153: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_153, data_out=>output_MAC_7_153);
	MAC_7_154: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_154, data_out=>output_MAC_7_154);
	MAC_7_155: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_155, data_out=>output_MAC_7_155);
	MAC_7_156: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_156, data_out=>output_MAC_7_156);
	MAC_7_157: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_157, data_out=>output_MAC_7_157);
	MAC_7_158: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_158, data_out=>output_MAC_7_158);
	MAC_7_159: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_159, data_out=>output_MAC_7_159);
	MAC_7_160: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_160, data_out=>output_MAC_7_160);
	MAC_7_161: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_161, data_out=>output_MAC_7_161);
	MAC_7_162: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_162, data_out=>output_MAC_7_162);
	MAC_7_163: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_163, data_out=>output_MAC_7_163);
	MAC_7_164: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_164, data_out=>output_MAC_7_164);
	MAC_7_165: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_165, data_out=>output_MAC_7_165);
	MAC_7_166: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_166, data_out=>output_MAC_7_166);
	MAC_7_167: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_167, data_out=>output_MAC_7_167);
	MAC_7_168: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_168, data_out=>output_MAC_7_168);
	MAC_7_169: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_169, data_out=>output_MAC_7_169);
	MAC_7_170: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_170, data_out=>output_MAC_7_170);
	MAC_7_171: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_171, data_out=>output_MAC_7_171);
	MAC_7_172: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_172, data_out=>output_MAC_7_172);
	MAC_7_173: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_173, data_out=>output_MAC_7_173);
	MAC_7_174: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_174, data_out=>output_MAC_7_174);
	MAC_7_175: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_175, data_out=>output_MAC_7_175);
	MAC_7_176: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_176, data_out=>output_MAC_7_176);
	MAC_7_177: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_177, data_out=>output_MAC_7_177);
	MAC_7_178: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_178, data_out=>output_MAC_7_178);
	MAC_7_179: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_179, data_out=>output_MAC_7_179);
	MAC_7_180: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_180, data_out=>output_MAC_7_180);
	MAC_7_181: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_181, data_out=>output_MAC_7_181);
	MAC_7_182: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_182, data_out=>output_MAC_7_182);
	MAC_7_183: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_183, data_out=>output_MAC_7_183);
	MAC_7_184: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_184, data_out=>output_MAC_7_184);
	MAC_7_185: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_185, data_out=>output_MAC_7_185);
	MAC_7_186: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_186, data_out=>output_MAC_7_186);
	MAC_7_187: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_187, data_out=>output_MAC_7_187);
	MAC_7_188: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_188, data_out=>output_MAC_7_188);
	MAC_7_189: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_189, data_out=>output_MAC_7_189);
	MAC_7_190: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_190, data_out=>output_MAC_7_190);
	MAC_7_191: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_191, data_out=>output_MAC_7_191);
	MAC_7_192: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_192, data_out=>output_MAC_7_192);
	MAC_7_193: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_193, data_out=>output_MAC_7_193);
	MAC_7_194: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_194, data_out=>output_MAC_7_194);
	MAC_7_195: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_195, data_out=>output_MAC_7_195);
	MAC_7_196: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_196, data_out=>output_MAC_7_196);
	MAC_7_197: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_197, data_out=>output_MAC_7_197);
	MAC_7_198: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_198, data_out=>output_MAC_7_198);
	MAC_7_199: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_199, data_out=>output_MAC_7_199);
	MAC_7_200: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_200, data_out=>output_MAC_7_200);
	MAC_7_201: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_201, data_out=>output_MAC_7_201);
	MAC_7_202: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_202, data_out=>output_MAC_7_202);
	MAC_7_203: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_203, data_out=>output_MAC_7_203);
	MAC_7_204: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_204, data_out=>output_MAC_7_204);
	MAC_7_205: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_205, data_out=>output_MAC_7_205);
	MAC_7_206: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_206, data_out=>output_MAC_7_206);
	MAC_7_207: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_207, data_out=>output_MAC_7_207);
	MAC_7_208: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_208, data_out=>output_MAC_7_208);
	MAC_7_209: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_209, data_out=>output_MAC_7_209);
	MAC_7_210: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_210, data_out=>output_MAC_7_210);
	MAC_7_211: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_211, data_out=>output_MAC_7_211);
	MAC_7_212: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_212, data_out=>output_MAC_7_212);
	MAC_7_213: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_213, data_out=>output_MAC_7_213);
	MAC_7_214: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_214, data_out=>output_MAC_7_214);
	MAC_7_215: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_215, data_out=>output_MAC_7_215);
	MAC_7_216: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_216, data_out=>output_MAC_7_216);
	MAC_7_217: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_217, data_out=>output_MAC_7_217);
	MAC_7_218: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_218, data_out=>output_MAC_7_218);
	MAC_7_219: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_219, data_out=>output_MAC_7_219);
	MAC_7_220: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_220, data_out=>output_MAC_7_220);
	MAC_7_221: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_221, data_out=>output_MAC_7_221);
	MAC_7_222: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_222, data_out=>output_MAC_7_222);
	MAC_7_223: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_223, data_out=>output_MAC_7_223);
	MAC_7_224: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_224, data_out=>output_MAC_7_224);
	MAC_7_225: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_225, data_out=>output_MAC_7_225);
	MAC_7_226: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_226, data_out=>output_MAC_7_226);
	MAC_7_227: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_227, data_out=>output_MAC_7_227);
	MAC_7_228: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_228, data_out=>output_MAC_7_228);
	MAC_7_229: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_229, data_out=>output_MAC_7_229);
	MAC_7_230: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_230, data_out=>output_MAC_7_230);
	MAC_7_231: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_231, data_out=>output_MAC_7_231);
	MAC_7_232: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_232, data_out=>output_MAC_7_232);
	MAC_7_233: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_233, data_out=>output_MAC_7_233);
	MAC_7_234: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_234, data_out=>output_MAC_7_234);
	MAC_7_235: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_235, data_out=>output_MAC_7_235);
	MAC_7_236: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_236, data_out=>output_MAC_7_236);
	MAC_7_237: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_237, data_out=>output_MAC_7_237);
	MAC_7_238: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_238, data_out=>output_MAC_7_238);
	MAC_7_239: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_239, data_out=>output_MAC_7_239);
	MAC_7_240: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_240, data_out=>output_MAC_7_240);
	MAC_7_241: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_241, data_out=>output_MAC_7_241);
	MAC_7_242: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_242, data_out=>output_MAC_7_242);
	MAC_7_243: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_243, data_out=>output_MAC_7_243);
	MAC_7_244: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_244, data_out=>output_MAC_7_244);
	MAC_7_245: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_245, data_out=>output_MAC_7_245);
	MAC_7_246: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_246, data_out=>output_MAC_7_246);
	MAC_7_247: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_247, data_out=>output_MAC_7_247);
	MAC_7_248: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_248, data_out=>output_MAC_7_248);
	MAC_7_249: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_249, data_out=>output_MAC_7_249);
	MAC_7_250: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_250, data_out=>output_MAC_7_250);
	MAC_7_251: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_251, data_out=>output_MAC_7_251);
	MAC_7_252: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_252, data_out=>output_MAC_7_252);
	MAC_7_253: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_253, data_out=>output_MAC_7_253);
	MAC_7_254: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_254, data_out=>output_MAC_7_254);
	MAC_7_255: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_255, data_out=>output_MAC_7_255);
	MAC_7_256: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_256, data_out=>output_MAC_7_256);
	MAC_7_257: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_257, data_out=>output_MAC_7_257);
	MAC_7_258: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_258, data_out=>output_MAC_7_258);
	MAC_7_259: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_259, data_out=>output_MAC_7_259);
	MAC_7_260: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_260, data_out=>output_MAC_7_260);
	MAC_7_261: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_261, data_out=>output_MAC_7_261);
	MAC_7_262: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_262, data_out=>output_MAC_7_262);
	MAC_7_263: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_263, data_out=>output_MAC_7_263);
	MAC_7_264: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_264, data_out=>output_MAC_7_264);
	MAC_7_265: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_265, data_out=>output_MAC_7_265);
	MAC_7_266: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_266, data_out=>output_MAC_7_266);
	MAC_7_267: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_267, data_out=>output_MAC_7_267);
	MAC_7_268: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_268, data_out=>output_MAC_7_268);
	MAC_7_269: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_269, data_out=>output_MAC_7_269);
	MAC_7_270: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_270, data_out=>output_MAC_7_270);
	MAC_7_271: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_271, data_out=>output_MAC_7_271);
	MAC_7_272: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_272, data_out=>output_MAC_7_272);
	MAC_7_273: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_273, data_out=>output_MAC_7_273);
	MAC_7_274: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_274, data_out=>output_MAC_7_274);
	MAC_7_275: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_275, data_out=>output_MAC_7_275);
	MAC_7_276: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_276, data_out=>output_MAC_7_276);
	MAC_7_277: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_277, data_out=>output_MAC_7_277);
	MAC_7_278: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_278, data_out=>output_MAC_7_278);
	MAC_7_279: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_279, data_out=>output_MAC_7_279);
	MAC_7_280: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_280, data_out=>output_MAC_7_280);
	MAC_7_281: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_281, data_out=>output_MAC_7_281);
	MAC_7_282: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_282, data_out=>output_MAC_7_282);
	MAC_7_283: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_283, data_out=>output_MAC_7_283);
	MAC_7_284: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_284, data_out=>output_MAC_7_284);
	MAC_7_285: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_285, data_out=>output_MAC_7_285);
	MAC_7_286: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_286, data_out=>output_MAC_7_286);
	MAC_7_287: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_287, data_out=>output_MAC_7_287);
	MAC_7_288: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_288, data_out=>output_MAC_7_288);
	MAC_7_289: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_289, data_out=>output_MAC_7_289);
	MAC_7_290: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_290, data_out=>output_MAC_7_290);
	MAC_7_291: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_291, data_out=>output_MAC_7_291);
	MAC_7_292: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_292, data_out=>output_MAC_7_292);
	MAC_7_293: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_293, data_out=>output_MAC_7_293);
	MAC_7_294: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_294, data_out=>output_MAC_7_294);
	MAC_7_295: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_295, data_out=>output_MAC_7_295);
	MAC_7_296: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_296, data_out=>output_MAC_7_296);
	MAC_7_297: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_297, data_out=>output_MAC_7_297);
	MAC_7_298: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_298, data_out=>output_MAC_7_298);
	MAC_7_299: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_299, data_out=>output_MAC_7_299);
	MAC_7_300: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_300, data_out=>output_MAC_7_300);
	MAC_7_301: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_301, data_out=>output_MAC_7_301);
	MAC_7_302: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_302, data_out=>output_MAC_7_302);
	MAC_7_303: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_303, data_out=>output_MAC_7_303);
	MAC_7_304: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_304, data_out=>output_MAC_7_304);
	MAC_7_305: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_305, data_out=>output_MAC_7_305);
	MAC_7_306: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_306, data_out=>output_MAC_7_306);
	MAC_7_307: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_307, data_out=>output_MAC_7_307);
	MAC_7_308: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_308, data_out=>output_MAC_7_308);
	MAC_7_309: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_309, data_out=>output_MAC_7_309);
	MAC_7_310: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_310, data_out=>output_MAC_7_310);
	MAC_7_311: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_311, data_out=>output_MAC_7_311);
	MAC_7_312: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_312, data_out=>output_MAC_7_312);
	MAC_7_313: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_313, data_out=>output_MAC_7_313);
	MAC_7_314: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_314, data_out=>output_MAC_7_314);
	MAC_7_315: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_315, data_out=>output_MAC_7_315);
	MAC_7_316: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_316, data_out=>output_MAC_7_316);
	MAC_7_317: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_317, data_out=>output_MAC_7_317);
	MAC_7_318: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_318, data_out=>output_MAC_7_318);
	MAC_7_319: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_319, data_out=>output_MAC_7_319);
	MAC_7_320: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_320, data_out=>output_MAC_7_320);
	MAC_7_321: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_321, data_out=>output_MAC_7_321);
	MAC_7_322: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_322, data_out=>output_MAC_7_322);
	MAC_7_323: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_323, data_out=>output_MAC_7_323);
	MAC_7_324: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_324, data_out=>output_MAC_7_324);
	MAC_7_325: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_325, data_out=>output_MAC_7_325);
	MAC_7_326: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_326, data_out=>output_MAC_7_326);
	MAC_7_327: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_327, data_out=>output_MAC_7_327);
	MAC_7_328: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_328, data_out=>output_MAC_7_328);
	MAC_7_329: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_329, data_out=>output_MAC_7_329);
	MAC_7_330: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_330, data_out=>output_MAC_7_330);
	MAC_7_331: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_331, data_out=>output_MAC_7_331);
	MAC_7_332: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_332, data_out=>output_MAC_7_332);
	MAC_7_333: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_333, data_out=>output_MAC_7_333);
	MAC_7_334: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_334, data_out=>output_MAC_7_334);
	MAC_7_335: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_335, data_out=>output_MAC_7_335);
	MAC_7_336: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_336, data_out=>output_MAC_7_336);
	MAC_7_337: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_337, data_out=>output_MAC_7_337);
	MAC_7_338: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_338, data_out=>output_MAC_7_338);
	MAC_7_339: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_339, data_out=>output_MAC_7_339);
	MAC_7_340: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_340, data_out=>output_MAC_7_340);
	MAC_7_341: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_341, data_out=>output_MAC_7_341);
	MAC_7_342: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_342, data_out=>output_MAC_7_342);
	MAC_7_343: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_343, data_out=>output_MAC_7_343);
	MAC_7_344: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_344, data_out=>output_MAC_7_344);
	MAC_7_345: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_345, data_out=>output_MAC_7_345);
	MAC_7_346: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_346, data_out=>output_MAC_7_346);
	MAC_7_347: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_347, data_out=>output_MAC_7_347);
	MAC_7_348: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_348, data_out=>output_MAC_7_348);
	MAC_7_349: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_349, data_out=>output_MAC_7_349);
	MAC_7_350: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_350, data_out=>output_MAC_7_350);
	MAC_7_351: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_351, data_out=>output_MAC_7_351);
	MAC_7_352: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_352, data_out=>output_MAC_7_352);
	MAC_7_353: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_353, data_out=>output_MAC_7_353);
	MAC_7_354: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_354, data_out=>output_MAC_7_354);
	MAC_7_355: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_355, data_out=>output_MAC_7_355);
	MAC_7_356: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_356, data_out=>output_MAC_7_356);
	MAC_7_357: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_357, data_out=>output_MAC_7_357);
	MAC_7_358: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_358, data_out=>output_MAC_7_358);
	MAC_7_359: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_359, data_out=>output_MAC_7_359);
	MAC_7_360: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_360, data_out=>output_MAC_7_360);
	MAC_7_361: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_361, data_out=>output_MAC_7_361);
	MAC_7_362: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_362, data_out=>output_MAC_7_362);
	MAC_7_363: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_363, data_out=>output_MAC_7_363);
	MAC_7_364: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_364, data_out=>output_MAC_7_364);
	MAC_7_365: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_365, data_out=>output_MAC_7_365);
	MAC_7_366: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_366, data_out=>output_MAC_7_366);
	MAC_7_367: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_367, data_out=>output_MAC_7_367);
	MAC_7_368: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_368, data_out=>output_MAC_7_368);
	MAC_7_369: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_369, data_out=>output_MAC_7_369);
	MAC_7_370: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_370, data_out=>output_MAC_7_370);
	MAC_7_371: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_371, data_out=>output_MAC_7_371);
	MAC_7_372: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_372, data_out=>output_MAC_7_372);
	MAC_7_373: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_373, data_out=>output_MAC_7_373);
	MAC_7_374: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_374, data_out=>output_MAC_7_374);
	MAC_7_375: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_375, data_out=>output_MAC_7_375);
	MAC_7_376: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_376, data_out=>output_MAC_7_376);
	MAC_7_377: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_377, data_out=>output_MAC_7_377);
	MAC_7_378: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_378, data_out=>output_MAC_7_378);
	MAC_7_379: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_379, data_out=>output_MAC_7_379);
	MAC_7_380: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_380, data_out=>output_MAC_7_380);
	MAC_7_381: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_381, data_out=>output_MAC_7_381);
	MAC_7_382: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_382, data_out=>output_MAC_7_382);
	MAC_7_383: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_383, data_out=>output_MAC_7_383);
	MAC_7_384: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_384, data_out=>output_MAC_7_384);
	MAC_7_385: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_385, data_out=>output_MAC_7_385);
	MAC_7_386: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_386, data_out=>output_MAC_7_386);
	MAC_7_387: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_387, data_out=>output_MAC_7_387);
	MAC_7_388: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_388, data_out=>output_MAC_7_388);
	MAC_7_389: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_389, data_out=>output_MAC_7_389);
	MAC_7_390: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_390, data_out=>output_MAC_7_390);
	MAC_7_391: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_391, data_out=>output_MAC_7_391);
	MAC_7_392: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_392, data_out=>output_MAC_7_392);
	MAC_7_393: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_393, data_out=>output_MAC_7_393);
	MAC_7_394: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_394, data_out=>output_MAC_7_394);
	MAC_7_395: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_395, data_out=>output_MAC_7_395);
	MAC_7_396: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_396, data_out=>output_MAC_7_396);
	MAC_7_397: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_397, data_out=>output_MAC_7_397);
	MAC_7_398: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_398, data_out=>output_MAC_7_398);
	MAC_7_399: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_399, data_out=>output_MAC_7_399);
	MAC_7_400: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_400, data_out=>output_MAC_7_400);
	MAC_7_401: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_401, data_out=>output_MAC_7_401);
	MAC_7_402: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_402, data_out=>output_MAC_7_402);
	MAC_7_403: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_403, data_out=>output_MAC_7_403);
	MAC_7_404: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_404, data_out=>output_MAC_7_404);
	MAC_7_405: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_405, data_out=>output_MAC_7_405);
	MAC_7_406: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_406, data_out=>output_MAC_7_406);
	MAC_7_407: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_407, data_out=>output_MAC_7_407);
	MAC_7_408: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_408, data_out=>output_MAC_7_408);
	MAC_7_409: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_409, data_out=>output_MAC_7_409);
	MAC_7_410: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_410, data_out=>output_MAC_7_410);
	MAC_7_411: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_411, data_out=>output_MAC_7_411);
	MAC_7_412: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_412, data_out=>output_MAC_7_412);
	MAC_7_413: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_413, data_out=>output_MAC_7_413);
	MAC_7_414: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_414, data_out=>output_MAC_7_414);
	MAC_7_415: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_415, data_out=>output_MAC_7_415);
	MAC_7_416: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_416, data_out=>output_MAC_7_416);
	MAC_7_417: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_417, data_out=>output_MAC_7_417);
	MAC_7_418: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_418, data_out=>output_MAC_7_418);
	MAC_7_419: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_419, data_out=>output_MAC_7_419);
	MAC_7_420: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_420, data_out=>output_MAC_7_420);
	MAC_7_421: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_421, data_out=>output_MAC_7_421);
	MAC_7_422: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_422, data_out=>output_MAC_7_422);
	MAC_7_423: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_423, data_out=>output_MAC_7_423);
	MAC_7_424: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_424, data_out=>output_MAC_7_424);
	MAC_7_425: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_425, data_out=>output_MAC_7_425);
	MAC_7_426: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_426, data_out=>output_MAC_7_426);
	MAC_7_427: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_427, data_out=>output_MAC_7_427);
	MAC_7_428: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_428, data_out=>output_MAC_7_428);
	MAC_7_429: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_429, data_out=>output_MAC_7_429);
	MAC_7_430: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_430, data_out=>output_MAC_7_430);
	MAC_7_431: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_431, data_out=>output_MAC_7_431);
	MAC_7_432: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_432, data_out=>output_MAC_7_432);
	MAC_7_433: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_433, data_out=>output_MAC_7_433);
	MAC_7_434: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_434, data_out=>output_MAC_7_434);
	MAC_7_435: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_435, data_out=>output_MAC_7_435);
	MAC_7_436: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_436, data_out=>output_MAC_7_436);
	MAC_7_437: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_437, data_out=>output_MAC_7_437);
	MAC_7_438: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_438, data_out=>output_MAC_7_438);
	MAC_7_439: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_439, data_out=>output_MAC_7_439);
	MAC_7_440: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_440, data_out=>output_MAC_7_440);
	MAC_7_441: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_441, data_out=>output_MAC_7_441);
	MAC_7_442: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_442, data_out=>output_MAC_7_442);
	MAC_7_443: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_443, data_out=>output_MAC_7_443);
	MAC_7_444: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_444, data_out=>output_MAC_7_444);
	MAC_7_445: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_445, data_out=>output_MAC_7_445);
	MAC_7_446: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_446, data_out=>output_MAC_7_446);
	MAC_7_447: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_447, data_out=>output_MAC_7_447);
	MAC_7_448: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_448, data_out=>output_MAC_7_448);
	MAC_7_449: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_449, data_out=>output_MAC_7_449);
	MAC_7_450: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_450, data_out=>output_MAC_7_450);
	MAC_7_451: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_451, data_out=>output_MAC_7_451);
	MAC_7_452: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_452, data_out=>output_MAC_7_452);
	MAC_7_453: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_453, data_out=>output_MAC_7_453);
	MAC_7_454: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_454, data_out=>output_MAC_7_454);
	MAC_7_455: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_455, data_out=>output_MAC_7_455);
	MAC_7_456: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_456, data_out=>output_MAC_7_456);
	MAC_7_457: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_457, data_out=>output_MAC_7_457);
	MAC_7_458: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_458, data_out=>output_MAC_7_458);
	MAC_7_459: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_459, data_out=>output_MAC_7_459);
	MAC_7_460: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_460, data_out=>output_MAC_7_460);
	MAC_7_461: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_461, data_out=>output_MAC_7_461);
	MAC_7_462: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_462, data_out=>output_MAC_7_462);
	MAC_7_463: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_463, data_out=>output_MAC_7_463);
	MAC_7_464: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_464, data_out=>output_MAC_7_464);
	MAC_7_465: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_465, data_out=>output_MAC_7_465);
	MAC_7_466: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_466, data_out=>output_MAC_7_466);
	MAC_7_467: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_467, data_out=>output_MAC_7_467);
	MAC_7_468: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_468, data_out=>output_MAC_7_468);
	MAC_7_469: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_469, data_out=>output_MAC_7_469);
	MAC_7_470: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_470, data_out=>output_MAC_7_470);
	MAC_7_471: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_471, data_out=>output_MAC_7_471);
	MAC_7_472: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_472, data_out=>output_MAC_7_472);
	MAC_7_473: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_473, data_out=>output_MAC_7_473);
	MAC_7_474: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_474, data_out=>output_MAC_7_474);
	MAC_7_475: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_475, data_out=>output_MAC_7_475);
	MAC_7_476: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_476, data_out=>output_MAC_7_476);
	MAC_7_477: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_477, data_out=>output_MAC_7_477);
	MAC_7_478: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_478, data_out=>output_MAC_7_478);
	MAC_7_479: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_479, data_out=>output_MAC_7_479);
	MAC_7_480: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_480, data_out=>output_MAC_7_480);
	MAC_7_481: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_481, data_out=>output_MAC_7_481);
	MAC_7_482: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_482, data_out=>output_MAC_7_482);
	MAC_7_483: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_483, data_out=>output_MAC_7_483);
	MAC_7_484: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_484, data_out=>output_MAC_7_484);
	MAC_7_485: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_485, data_out=>output_MAC_7_485);
	MAC_7_486: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_486, data_out=>output_MAC_7_486);
	MAC_7_487: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_487, data_out=>output_MAC_7_487);
	MAC_7_488: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_488, data_out=>output_MAC_7_488);
	MAC_7_489: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_489, data_out=>output_MAC_7_489);
	MAC_7_490: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_490, data_out=>output_MAC_7_490);
	MAC_7_491: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_491, data_out=>output_MAC_7_491);
	MAC_7_492: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_492, data_out=>output_MAC_7_492);
	MAC_7_493: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_493, data_out=>output_MAC_7_493);
	MAC_7_494: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_494, data_out=>output_MAC_7_494);
	MAC_7_495: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_495, data_out=>output_MAC_7_495);
	MAC_7_496: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_496, data_out=>output_MAC_7_496);
	MAC_7_497: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_497, data_out=>output_MAC_7_497);
	MAC_7_498: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_498, data_out=>output_MAC_7_498);
	MAC_7_499: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_499, data_out=>output_MAC_7_499);
	MAC_7_500: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_500, data_out=>output_MAC_7_500);
	MAC_7_501: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_501, data_out=>output_MAC_7_501);
	MAC_7_502: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_502, data_out=>output_MAC_7_502);
	MAC_7_503: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_503, data_out=>output_MAC_7_503);
	MAC_7_504: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_504, data_out=>output_MAC_7_504);
	MAC_7_505: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_505, data_out=>output_MAC_7_505);
	MAC_7_506: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_506, data_out=>output_MAC_7_506);
	MAC_7_507: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_507, data_out=>output_MAC_7_507);
	MAC_7_508: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_508, data_out=>output_MAC_7_508);
	MAC_7_509: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_509, data_out=>output_MAC_7_509);
	MAC_7_510: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_510, data_out=>output_MAC_7_510);
	MAC_7_511: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_511, data_out=>output_MAC_7_511);
	MAC_7_512: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_512, data_out=>output_MAC_7_512);
	MAC_7_513: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_513, data_out=>output_MAC_7_513);
	MAC_7_514: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_514, data_out=>output_MAC_7_514);
	MAC_7_515: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_515, data_out=>output_MAC_7_515);
	MAC_7_516: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_516, data_out=>output_MAC_7_516);
	MAC_7_517: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_517, data_out=>output_MAC_7_517);
	MAC_7_518: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_518, data_out=>output_MAC_7_518);
	MAC_7_519: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_519, data_out=>output_MAC_7_519);
	MAC_7_520: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_520, data_out=>output_MAC_7_520);
	MAC_7_521: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_521, data_out=>output_MAC_7_521);
	MAC_7_522: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_522, data_out=>output_MAC_7_522);
	MAC_7_523: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_523, data_out=>output_MAC_7_523);
	MAC_7_524: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_524, data_out=>output_MAC_7_524);
	MAC_7_525: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_525, data_out=>output_MAC_7_525);
	MAC_7_526: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_526, data_out=>output_MAC_7_526);
	MAC_7_527: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_527, data_out=>output_MAC_7_527);
	MAC_7_528: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_528, data_out=>output_MAC_7_528);
	MAC_7_529: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_529, data_out=>output_MAC_7_529);
	MAC_7_530: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_530, data_out=>output_MAC_7_530);
	MAC_7_531: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_531, data_out=>output_MAC_7_531);
	MAC_7_532: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_532, data_out=>output_MAC_7_532);
	MAC_7_533: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_533, data_out=>output_MAC_7_533);
	MAC_7_534: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_534, data_out=>output_MAC_7_534);
	MAC_7_535: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_535, data_out=>output_MAC_7_535);
	MAC_7_536: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_536, data_out=>output_MAC_7_536);
	MAC_7_537: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_537, data_out=>output_MAC_7_537);
	MAC_7_538: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_538, data_out=>output_MAC_7_538);
	MAC_7_539: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_539, data_out=>output_MAC_7_539);
	MAC_7_540: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_540, data_out=>output_MAC_7_540);
	MAC_7_541: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_541, data_out=>output_MAC_7_541);
	MAC_7_542: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_542, data_out=>output_MAC_7_542);
	MAC_7_543: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_543, data_out=>output_MAC_7_543);
	MAC_7_544: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_544, data_out=>output_MAC_7_544);
	MAC_7_545: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_545, data_out=>output_MAC_7_545);
	MAC_7_546: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_546, data_out=>output_MAC_7_546);
	MAC_7_547: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_547, data_out=>output_MAC_7_547);
	MAC_7_548: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_548, data_out=>output_MAC_7_548);
	MAC_7_549: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_549, data_out=>output_MAC_7_549);
	MAC_7_550: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_550, data_out=>output_MAC_7_550);
	MAC_7_551: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_551, data_out=>output_MAC_7_551);
	MAC_7_552: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_552, data_out=>output_MAC_7_552);
	MAC_7_553: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_553, data_out=>output_MAC_7_553);
	MAC_7_554: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_554, data_out=>output_MAC_7_554);
	MAC_7_555: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_555, data_out=>output_MAC_7_555);
	MAC_7_556: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_556, data_out=>output_MAC_7_556);
	MAC_7_557: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_557, data_out=>output_MAC_7_557);
	MAC_7_558: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_558, data_out=>output_MAC_7_558);
	MAC_7_559: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_559, data_out=>output_MAC_7_559);
	MAC_7_560: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_560, data_out=>output_MAC_7_560);
	MAC_7_561: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_561, data_out=>output_MAC_7_561);
	MAC_7_562: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_562, data_out=>output_MAC_7_562);
	MAC_7_563: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_563, data_out=>output_MAC_7_563);
	MAC_7_564: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_564, data_out=>output_MAC_7_564);
	MAC_7_565: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_565, data_out=>output_MAC_7_565);
	MAC_7_566: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_566, data_out=>output_MAC_7_566);
	MAC_7_567: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_567, data_out=>output_MAC_7_567);
	MAC_7_568: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_568, data_out=>output_MAC_7_568);
	MAC_7_569: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_569, data_out=>output_MAC_7_569);
	MAC_7_570: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_570, data_out=>output_MAC_7_570);
	MAC_7_571: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_571, data_out=>output_MAC_7_571);
	MAC_7_572: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_572, data_out=>output_MAC_7_572);
	MAC_7_573: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_573, data_out=>output_MAC_7_573);
	MAC_7_574: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_574, data_out=>output_MAC_7_574);
	MAC_7_575: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_575, data_out=>output_MAC_7_575);
	MAC_7_576: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_576, data_out=>output_MAC_7_576);
	MAC_7_577: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_577, data_out=>output_MAC_7_577);
	MAC_7_578: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_578, data_out=>output_MAC_7_578);
	MAC_7_579: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_579, data_out=>output_MAC_7_579);
	MAC_7_580: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_580, data_out=>output_MAC_7_580);
	MAC_7_581: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_581, data_out=>output_MAC_7_581);
	MAC_7_582: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_582, data_out=>output_MAC_7_582);
	MAC_7_583: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_583, data_out=>output_MAC_7_583);
	MAC_7_584: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_584, data_out=>output_MAC_7_584);
	MAC_7_585: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_585, data_out=>output_MAC_7_585);
	MAC_7_586: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_586, data_out=>output_MAC_7_586);
	MAC_7_587: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_587, data_out=>output_MAC_7_587);
	MAC_7_588: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_588, data_out=>output_MAC_7_588);
	MAC_7_589: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_589, data_out=>output_MAC_7_589);
	MAC_7_590: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_590, data_out=>output_MAC_7_590);
	MAC_7_591: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_591, data_out=>output_MAC_7_591);
	MAC_7_592: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_592, data_out=>output_MAC_7_592);
	MAC_7_593: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_593, data_out=>output_MAC_7_593);
	MAC_7_594: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_594, data_out=>output_MAC_7_594);
	MAC_7_595: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_595, data_out=>output_MAC_7_595);
	MAC_7_596: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_596, data_out=>output_MAC_7_596);
	MAC_7_597: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_597, data_out=>output_MAC_7_597);
	MAC_7_598: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_598, data_out=>output_MAC_7_598);
	MAC_7_599: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_599, data_out=>output_MAC_7_599);
	MAC_7_600: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_600, data_out=>output_MAC_7_600);
	MAC_7_601: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_601, data_out=>output_MAC_7_601);
	MAC_7_602: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_602, data_out=>output_MAC_7_602);
	MAC_7_603: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_603, data_out=>output_MAC_7_603);
	MAC_7_604: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_604, data_out=>output_MAC_7_604);
	MAC_7_605: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_605, data_out=>output_MAC_7_605);
	MAC_7_606: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_606, data_out=>output_MAC_7_606);
	MAC_7_607: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_607, data_out=>output_MAC_7_607);
	MAC_7_608: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_608, data_out=>output_MAC_7_608);
	MAC_7_609: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_609, data_out=>output_MAC_7_609);
	MAC_7_610: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_610, data_out=>output_MAC_7_610);
	MAC_7_611: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_611, data_out=>output_MAC_7_611);
	MAC_7_612: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_612, data_out=>output_MAC_7_612);
	MAC_7_613: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_613, data_out=>output_MAC_7_613);
	MAC_7_614: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_614, data_out=>output_MAC_7_614);
	MAC_7_615: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_615, data_out=>output_MAC_7_615);
	MAC_7_616: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_616, data_out=>output_MAC_7_616);
	MAC_7_617: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_617, data_out=>output_MAC_7_617);
	MAC_7_618: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_618, data_out=>output_MAC_7_618);
	MAC_7_619: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_619, data_out=>output_MAC_7_619);
	MAC_7_620: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_620, data_out=>output_MAC_7_620);
	MAC_7_621: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_621, data_out=>output_MAC_7_621);
	MAC_7_622: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_622, data_out=>output_MAC_7_622);
	MAC_7_623: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_623, data_out=>output_MAC_7_623);
	MAC_7_624: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_624, data_out=>output_MAC_7_624);
	MAC_7_625: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_625, data_out=>output_MAC_7_625);
	MAC_7_626: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_626, data_out=>output_MAC_7_626);
	MAC_7_627: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_627, data_out=>output_MAC_7_627);
	MAC_7_628: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_628, data_out=>output_MAC_7_628);
	MAC_7_629: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_629, data_out=>output_MAC_7_629);
	MAC_7_630: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_630, data_out=>output_MAC_7_630);
	MAC_7_631: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_631, data_out=>output_MAC_7_631);
	MAC_7_632: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_632, data_out=>output_MAC_7_632);
	MAC_7_633: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_633, data_out=>output_MAC_7_633);
	MAC_7_634: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_634, data_out=>output_MAC_7_634);
	MAC_7_635: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_635, data_out=>output_MAC_7_635);
	MAC_7_636: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_636, data_out=>output_MAC_7_636);
	MAC_7_637: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_637, data_out=>output_MAC_7_637);
	MAC_7_638: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_638, data_out=>output_MAC_7_638);
	MAC_7_639: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_639, data_out=>output_MAC_7_639);
	MAC_7_640: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_640, data_out=>output_MAC_7_640);
	MAC_7_641: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_641, data_out=>output_MAC_7_641);
	MAC_7_642: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_642, data_out=>output_MAC_7_642);
	MAC_7_643: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_643, data_out=>output_MAC_7_643);
	MAC_7_644: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_644, data_out=>output_MAC_7_644);
	MAC_7_645: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_645, data_out=>output_MAC_7_645);
	MAC_7_646: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_646, data_out=>output_MAC_7_646);
	MAC_7_647: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_647, data_out=>output_MAC_7_647);
	MAC_7_648: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_648, data_out=>output_MAC_7_648);
	MAC_7_649: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_649, data_out=>output_MAC_7_649);
	MAC_7_650: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_650, data_out=>output_MAC_7_650);
	MAC_7_651: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_651, data_out=>output_MAC_7_651);
	MAC_7_652: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_652, data_out=>output_MAC_7_652);
	MAC_7_653: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_653, data_out=>output_MAC_7_653);
	MAC_7_654: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_654, data_out=>output_MAC_7_654);
	MAC_7_655: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_655, data_out=>output_MAC_7_655);
	MAC_7_656: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_656, data_out=>output_MAC_7_656);
	MAC_7_657: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_657, data_out=>output_MAC_7_657);
	MAC_7_658: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_658, data_out=>output_MAC_7_658);
	MAC_7_659: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_659, data_out=>output_MAC_7_659);
	MAC_7_660: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_660, data_out=>output_MAC_7_660);
	MAC_7_661: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_661, data_out=>output_MAC_7_661);
	MAC_7_662: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_662, data_out=>output_MAC_7_662);
	MAC_7_663: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_663, data_out=>output_MAC_7_663);
	MAC_7_664: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_664, data_out=>output_MAC_7_664);
	MAC_7_665: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_665, data_out=>output_MAC_7_665);
	MAC_7_666: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_666, data_out=>output_MAC_7_666);
	MAC_7_667: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_667, data_out=>output_MAC_7_667);
	MAC_7_668: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_668, data_out=>output_MAC_7_668);
	MAC_7_669: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_669, data_out=>output_MAC_7_669);
	MAC_7_670: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_670, data_out=>output_MAC_7_670);
	MAC_7_671: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_671, data_out=>output_MAC_7_671);
	MAC_7_672: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_672, data_out=>output_MAC_7_672);
	MAC_7_673: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_673, data_out=>output_MAC_7_673);
	MAC_7_674: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_674, data_out=>output_MAC_7_674);
	MAC_7_675: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_675, data_out=>output_MAC_7_675);
	MAC_7_676: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_676, data_out=>output_MAC_7_676);
	MAC_7_677: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_677, data_out=>output_MAC_7_677);
	MAC_7_678: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_678, data_out=>output_MAC_7_678);
	MAC_7_679: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_679, data_out=>output_MAC_7_679);
	MAC_7_680: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_680, data_out=>output_MAC_7_680);
	MAC_7_681: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_681, data_out=>output_MAC_7_681);
	MAC_7_682: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_682, data_out=>output_MAC_7_682);
	MAC_7_683: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_683, data_out=>output_MAC_7_683);
	MAC_7_684: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_684, data_out=>output_MAC_7_684);
	MAC_7_685: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_685, data_out=>output_MAC_7_685);
	MAC_7_686: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_686, data_out=>output_MAC_7_686);
	MAC_7_687: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_687, data_out=>output_MAC_7_687);
	MAC_7_688: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_688, data_out=>output_MAC_7_688);
	MAC_7_689: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_689, data_out=>output_MAC_7_689);
	MAC_7_690: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_690, data_out=>output_MAC_7_690);
	MAC_7_691: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_691, data_out=>output_MAC_7_691);
	MAC_7_692: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_692, data_out=>output_MAC_7_692);
	MAC_7_693: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_693, data_out=>output_MAC_7_693);
	MAC_7_694: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_694, data_out=>output_MAC_7_694);
	MAC_7_695: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_695, data_out=>output_MAC_7_695);
	MAC_7_696: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_696, data_out=>output_MAC_7_696);
	MAC_7_697: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_697, data_out=>output_MAC_7_697);
	MAC_7_698: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_698, data_out=>output_MAC_7_698);
	MAC_7_699: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_699, data_out=>output_MAC_7_699);
	MAC_7_700: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_700, data_out=>output_MAC_7_700);
	MAC_7_701: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_701, data_out=>output_MAC_7_701);
	MAC_7_702: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_702, data_out=>output_MAC_7_702);
	MAC_7_703: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_703, data_out=>output_MAC_7_703);
	MAC_7_704: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_704, data_out=>output_MAC_7_704);
	MAC_7_705: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_705, data_out=>output_MAC_7_705);
	MAC_7_706: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_706, data_out=>output_MAC_7_706);
	MAC_7_707: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_707, data_out=>output_MAC_7_707);
	MAC_7_708: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_708, data_out=>output_MAC_7_708);
	MAC_7_709: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_709, data_out=>output_MAC_7_709);
	MAC_7_710: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_710, data_out=>output_MAC_7_710);
	MAC_7_711: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_711, data_out=>output_MAC_7_711);
	MAC_7_712: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_712, data_out=>output_MAC_7_712);
	MAC_7_713: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_713, data_out=>output_MAC_7_713);
	MAC_7_714: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_714, data_out=>output_MAC_7_714);
	MAC_7_715: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_715, data_out=>output_MAC_7_715);
	MAC_7_716: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_716, data_out=>output_MAC_7_716);
	MAC_7_717: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_717, data_out=>output_MAC_7_717);
	MAC_7_718: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_718, data_out=>output_MAC_7_718);
	MAC_7_719: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_719, data_out=>output_MAC_7_719);
	MAC_7_720: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_720, data_out=>output_MAC_7_720);
	MAC_7_721: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_721, data_out=>output_MAC_7_721);
	MAC_7_722: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_722, data_out=>output_MAC_7_722);
	MAC_7_723: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_723, data_out=>output_MAC_7_723);
	MAC_7_724: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_724, data_out=>output_MAC_7_724);
	MAC_7_725: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_725, data_out=>output_MAC_7_725);
	MAC_7_726: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_726, data_out=>output_MAC_7_726);
	MAC_7_727: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_727, data_out=>output_MAC_7_727);
	MAC_7_728: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_728, data_out=>output_MAC_7_728);
	MAC_7_729: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_729, data_out=>output_MAC_7_729);
	MAC_7_730: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_730, data_out=>output_MAC_7_730);
	MAC_7_731: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_731, data_out=>output_MAC_7_731);
	MAC_7_732: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_732, data_out=>output_MAC_7_732);
	MAC_7_733: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_733, data_out=>output_MAC_7_733);
	MAC_7_734: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_734, data_out=>output_MAC_7_734);
	MAC_7_735: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_735, data_out=>output_MAC_7_735);
	MAC_7_736: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_736, data_out=>output_MAC_7_736);
	MAC_7_737: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_737, data_out=>output_MAC_7_737);
	MAC_7_738: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_738, data_out=>output_MAC_7_738);
	MAC_7_739: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_739, data_out=>output_MAC_7_739);
	MAC_7_740: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_740, data_out=>output_MAC_7_740);
	MAC_7_741: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_741, data_out=>output_MAC_7_741);
	MAC_7_742: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_742, data_out=>output_MAC_7_742);
	MAC_7_743: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_743, data_out=>output_MAC_7_743);
	MAC_7_744: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_744, data_out=>output_MAC_7_744);
	MAC_7_745: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_745, data_out=>output_MAC_7_745);
	MAC_7_746: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_746, data_out=>output_MAC_7_746);
	MAC_7_747: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_747, data_out=>output_MAC_7_747);
	MAC_7_748: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_748, data_out=>output_MAC_7_748);
	MAC_7_749: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_749, data_out=>output_MAC_7_749);
	MAC_7_750: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_750, data_out=>output_MAC_7_750);
	MAC_7_751: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_751, data_out=>output_MAC_7_751);
	MAC_7_752: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_752, data_out=>output_MAC_7_752);
	MAC_7_753: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_753, data_out=>output_MAC_7_753);
	MAC_7_754: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_754, data_out=>output_MAC_7_754);
	MAC_7_755: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_755, data_out=>output_MAC_7_755);
	MAC_7_756: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_756, data_out=>output_MAC_7_756);
	MAC_7_757: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_757, data_out=>output_MAC_7_757);
	MAC_7_758: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_758, data_out=>output_MAC_7_758);
	MAC_7_759: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_759, data_out=>output_MAC_7_759);
	MAC_7_760: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_760, data_out=>output_MAC_7_760);
	MAC_7_761: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_761, data_out=>output_MAC_7_761);
	MAC_7_762: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_762, data_out=>output_MAC_7_762);
	MAC_7_763: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_763, data_out=>output_MAC_7_763);
	MAC_7_764: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_764, data_out=>output_MAC_7_764);
	MAC_7_765: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_765, data_out=>output_MAC_7_765);
	MAC_7_766: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_766, data_out=>output_MAC_7_766);
	MAC_7_767: MAC GENERIC MAP(data_size=>8, acc_size=>32)
			PORT MAP(CLK=>CLK, RST_n=>RST_n, ENABLE=>ENABLE, data_in_A=>input_row_7, data_in_B=>input_col_767, data_out=>output_MAC_7_767);

	mux_row_0: mux_768to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_0_0, I1=>output_MAC_0_1, I2=>output_MAC_0_2, I3=>output_MAC_0_3, I4=>output_MAC_0_4, I5=>output_MAC_0_5, I6=>output_MAC_0_6, I7=>output_MAC_0_7, I8=>output_MAC_0_8, I9=>output_MAC_0_9, I10=>output_MAC_0_10, I11=>output_MAC_0_11, I12=>output_MAC_0_12, I13=>output_MAC_0_13, I14=>output_MAC_0_14, I15=>output_MAC_0_15, I16=>output_MAC_0_16, I17=>output_MAC_0_17, I18=>output_MAC_0_18, I19=>output_MAC_0_19, I20=>output_MAC_0_20, I21=>output_MAC_0_21, I22=>output_MAC_0_22, I23=>output_MAC_0_23, I24=>output_MAC_0_24, I25=>output_MAC_0_25, I26=>output_MAC_0_26, I27=>output_MAC_0_27, I28=>output_MAC_0_28, I29=>output_MAC_0_29, I30=>output_MAC_0_30, I31=>output_MAC_0_31, I32=>output_MAC_0_32, I33=>output_MAC_0_33, I34=>output_MAC_0_34, I35=>output_MAC_0_35, I36=>output_MAC_0_36, I37=>output_MAC_0_37, I38=>output_MAC_0_38, I39=>output_MAC_0_39, I40=>output_MAC_0_40, I41=>output_MAC_0_41, I42=>output_MAC_0_42, I43=>output_MAC_0_43, I44=>output_MAC_0_44, I45=>output_MAC_0_45, I46=>output_MAC_0_46, I47=>output_MAC_0_47, I48=>output_MAC_0_48, I49=>output_MAC_0_49, I50=>output_MAC_0_50, I51=>output_MAC_0_51, I52=>output_MAC_0_52, I53=>output_MAC_0_53, I54=>output_MAC_0_54, I55=>output_MAC_0_55, I56=>output_MAC_0_56, I57=>output_MAC_0_57, I58=>output_MAC_0_58, I59=>output_MAC_0_59, I60=>output_MAC_0_60, I61=>output_MAC_0_61, I62=>output_MAC_0_62, I63=>output_MAC_0_63, I64=>output_MAC_0_64, I65=>output_MAC_0_65, I66=>output_MAC_0_66, I67=>output_MAC_0_67, I68=>output_MAC_0_68, I69=>output_MAC_0_69, I70=>output_MAC_0_70, I71=>output_MAC_0_71, I72=>output_MAC_0_72, I73=>output_MAC_0_73, I74=>output_MAC_0_74, I75=>output_MAC_0_75, I76=>output_MAC_0_76, I77=>output_MAC_0_77, I78=>output_MAC_0_78, I79=>output_MAC_0_79, I80=>output_MAC_0_80, I81=>output_MAC_0_81, I82=>output_MAC_0_82, I83=>output_MAC_0_83, I84=>output_MAC_0_84, I85=>output_MAC_0_85, I86=>output_MAC_0_86, I87=>output_MAC_0_87, I88=>output_MAC_0_88, I89=>output_MAC_0_89, I90=>output_MAC_0_90, I91=>output_MAC_0_91, I92=>output_MAC_0_92, I93=>output_MAC_0_93, I94=>output_MAC_0_94, I95=>output_MAC_0_95, I96=>output_MAC_0_96, I97=>output_MAC_0_97, I98=>output_MAC_0_98, I99=>output_MAC_0_99, I100=>output_MAC_0_100, I101=>output_MAC_0_101, I102=>output_MAC_0_102, I103=>output_MAC_0_103, I104=>output_MAC_0_104, I105=>output_MAC_0_105, I106=>output_MAC_0_106, I107=>output_MAC_0_107, I108=>output_MAC_0_108, I109=>output_MAC_0_109, I110=>output_MAC_0_110, I111=>output_MAC_0_111, I112=>output_MAC_0_112, I113=>output_MAC_0_113, I114=>output_MAC_0_114, I115=>output_MAC_0_115, I116=>output_MAC_0_116, I117=>output_MAC_0_117, I118=>output_MAC_0_118, I119=>output_MAC_0_119, I120=>output_MAC_0_120, I121=>output_MAC_0_121, I122=>output_MAC_0_122, I123=>output_MAC_0_123, I124=>output_MAC_0_124, I125=>output_MAC_0_125, I126=>output_MAC_0_126, I127=>output_MAC_0_127, I128=>output_MAC_0_128, I129=>output_MAC_0_129, I130=>output_MAC_0_130, I131=>output_MAC_0_131, I132=>output_MAC_0_132, I133=>output_MAC_0_133, I134=>output_MAC_0_134, I135=>output_MAC_0_135, I136=>output_MAC_0_136, I137=>output_MAC_0_137, I138=>output_MAC_0_138, I139=>output_MAC_0_139, I140=>output_MAC_0_140, I141=>output_MAC_0_141, I142=>output_MAC_0_142, I143=>output_MAC_0_143, I144=>output_MAC_0_144, I145=>output_MAC_0_145, I146=>output_MAC_0_146, I147=>output_MAC_0_147, I148=>output_MAC_0_148, I149=>output_MAC_0_149, I150=>output_MAC_0_150, I151=>output_MAC_0_151, I152=>output_MAC_0_152, I153=>output_MAC_0_153, I154=>output_MAC_0_154, I155=>output_MAC_0_155, I156=>output_MAC_0_156, I157=>output_MAC_0_157, I158=>output_MAC_0_158, I159=>output_MAC_0_159, I160=>output_MAC_0_160, I161=>output_MAC_0_161, I162=>output_MAC_0_162, I163=>output_MAC_0_163, I164=>output_MAC_0_164, I165=>output_MAC_0_165, I166=>output_MAC_0_166, I167=>output_MAC_0_167, I168=>output_MAC_0_168, I169=>output_MAC_0_169, I170=>output_MAC_0_170, I171=>output_MAC_0_171, I172=>output_MAC_0_172, I173=>output_MAC_0_173, I174=>output_MAC_0_174, I175=>output_MAC_0_175, I176=>output_MAC_0_176, I177=>output_MAC_0_177, I178=>output_MAC_0_178, I179=>output_MAC_0_179, I180=>output_MAC_0_180, I181=>output_MAC_0_181, I182=>output_MAC_0_182, I183=>output_MAC_0_183, I184=>output_MAC_0_184, I185=>output_MAC_0_185, I186=>output_MAC_0_186, I187=>output_MAC_0_187, I188=>output_MAC_0_188, I189=>output_MAC_0_189, I190=>output_MAC_0_190, I191=>output_MAC_0_191, I192=>output_MAC_0_192, I193=>output_MAC_0_193, I194=>output_MAC_0_194, I195=>output_MAC_0_195, I196=>output_MAC_0_196, I197=>output_MAC_0_197, I198=>output_MAC_0_198, I199=>output_MAC_0_199, I200=>output_MAC_0_200, I201=>output_MAC_0_201, I202=>output_MAC_0_202, I203=>output_MAC_0_203, I204=>output_MAC_0_204, I205=>output_MAC_0_205, I206=>output_MAC_0_206, I207=>output_MAC_0_207, I208=>output_MAC_0_208, I209=>output_MAC_0_209, I210=>output_MAC_0_210, I211=>output_MAC_0_211, I212=>output_MAC_0_212, I213=>output_MAC_0_213, I214=>output_MAC_0_214, I215=>output_MAC_0_215, I216=>output_MAC_0_216, I217=>output_MAC_0_217, I218=>output_MAC_0_218, I219=>output_MAC_0_219, I220=>output_MAC_0_220, I221=>output_MAC_0_221, I222=>output_MAC_0_222, I223=>output_MAC_0_223, I224=>output_MAC_0_224, I225=>output_MAC_0_225, I226=>output_MAC_0_226, I227=>output_MAC_0_227, I228=>output_MAC_0_228, I229=>output_MAC_0_229, I230=>output_MAC_0_230, I231=>output_MAC_0_231, I232=>output_MAC_0_232, I233=>output_MAC_0_233, I234=>output_MAC_0_234, I235=>output_MAC_0_235, I236=>output_MAC_0_236, I237=>output_MAC_0_237, I238=>output_MAC_0_238, I239=>output_MAC_0_239, I240=>output_MAC_0_240, I241=>output_MAC_0_241, I242=>output_MAC_0_242, I243=>output_MAC_0_243, I244=>output_MAC_0_244, I245=>output_MAC_0_245, I246=>output_MAC_0_246, I247=>output_MAC_0_247, I248=>output_MAC_0_248, I249=>output_MAC_0_249, I250=>output_MAC_0_250, I251=>output_MAC_0_251, I252=>output_MAC_0_252, I253=>output_MAC_0_253, I254=>output_MAC_0_254, I255=>output_MAC_0_255, I256=>output_MAC_0_256, I257=>output_MAC_0_257, I258=>output_MAC_0_258, I259=>output_MAC_0_259, I260=>output_MAC_0_260, I261=>output_MAC_0_261, I262=>output_MAC_0_262, I263=>output_MAC_0_263, I264=>output_MAC_0_264, I265=>output_MAC_0_265, I266=>output_MAC_0_266, I267=>output_MAC_0_267, I268=>output_MAC_0_268, I269=>output_MAC_0_269, I270=>output_MAC_0_270, I271=>output_MAC_0_271, I272=>output_MAC_0_272, I273=>output_MAC_0_273, I274=>output_MAC_0_274, I275=>output_MAC_0_275, I276=>output_MAC_0_276, I277=>output_MAC_0_277, I278=>output_MAC_0_278, I279=>output_MAC_0_279, I280=>output_MAC_0_280, I281=>output_MAC_0_281, I282=>output_MAC_0_282, I283=>output_MAC_0_283, I284=>output_MAC_0_284, I285=>output_MAC_0_285, I286=>output_MAC_0_286, I287=>output_MAC_0_287, I288=>output_MAC_0_288, I289=>output_MAC_0_289, I290=>output_MAC_0_290, I291=>output_MAC_0_291, I292=>output_MAC_0_292, I293=>output_MAC_0_293, I294=>output_MAC_0_294, I295=>output_MAC_0_295, I296=>output_MAC_0_296, I297=>output_MAC_0_297, I298=>output_MAC_0_298, I299=>output_MAC_0_299, I300=>output_MAC_0_300, I301=>output_MAC_0_301, I302=>output_MAC_0_302, I303=>output_MAC_0_303, I304=>output_MAC_0_304, I305=>output_MAC_0_305, I306=>output_MAC_0_306, I307=>output_MAC_0_307, I308=>output_MAC_0_308, I309=>output_MAC_0_309, I310=>output_MAC_0_310, I311=>output_MAC_0_311, I312=>output_MAC_0_312, I313=>output_MAC_0_313, I314=>output_MAC_0_314, I315=>output_MAC_0_315, I316=>output_MAC_0_316, I317=>output_MAC_0_317, I318=>output_MAC_0_318, I319=>output_MAC_0_319, I320=>output_MAC_0_320, I321=>output_MAC_0_321, I322=>output_MAC_0_322, I323=>output_MAC_0_323, I324=>output_MAC_0_324, I325=>output_MAC_0_325, I326=>output_MAC_0_326, I327=>output_MAC_0_327, I328=>output_MAC_0_328, I329=>output_MAC_0_329, I330=>output_MAC_0_330, I331=>output_MAC_0_331, I332=>output_MAC_0_332, I333=>output_MAC_0_333, I334=>output_MAC_0_334, I335=>output_MAC_0_335, I336=>output_MAC_0_336, I337=>output_MAC_0_337, I338=>output_MAC_0_338, I339=>output_MAC_0_339, I340=>output_MAC_0_340, I341=>output_MAC_0_341, I342=>output_MAC_0_342, I343=>output_MAC_0_343, I344=>output_MAC_0_344, I345=>output_MAC_0_345, I346=>output_MAC_0_346, I347=>output_MAC_0_347, I348=>output_MAC_0_348, I349=>output_MAC_0_349, I350=>output_MAC_0_350, I351=>output_MAC_0_351, I352=>output_MAC_0_352, I353=>output_MAC_0_353, I354=>output_MAC_0_354, I355=>output_MAC_0_355, I356=>output_MAC_0_356, I357=>output_MAC_0_357, I358=>output_MAC_0_358, I359=>output_MAC_0_359, I360=>output_MAC_0_360, I361=>output_MAC_0_361, I362=>output_MAC_0_362, I363=>output_MAC_0_363, I364=>output_MAC_0_364, I365=>output_MAC_0_365, I366=>output_MAC_0_366, I367=>output_MAC_0_367, I368=>output_MAC_0_368, I369=>output_MAC_0_369, I370=>output_MAC_0_370, I371=>output_MAC_0_371, I372=>output_MAC_0_372, I373=>output_MAC_0_373, I374=>output_MAC_0_374, I375=>output_MAC_0_375, I376=>output_MAC_0_376, I377=>output_MAC_0_377, I378=>output_MAC_0_378, I379=>output_MAC_0_379, I380=>output_MAC_0_380, I381=>output_MAC_0_381, I382=>output_MAC_0_382, I383=>output_MAC_0_383, I384=>output_MAC_0_384, I385=>output_MAC_0_385, I386=>output_MAC_0_386, I387=>output_MAC_0_387, I388=>output_MAC_0_388, I389=>output_MAC_0_389, I390=>output_MAC_0_390, I391=>output_MAC_0_391, I392=>output_MAC_0_392, I393=>output_MAC_0_393, I394=>output_MAC_0_394, I395=>output_MAC_0_395, I396=>output_MAC_0_396, I397=>output_MAC_0_397, I398=>output_MAC_0_398, I399=>output_MAC_0_399, I400=>output_MAC_0_400, I401=>output_MAC_0_401, I402=>output_MAC_0_402, I403=>output_MAC_0_403, I404=>output_MAC_0_404, I405=>output_MAC_0_405, I406=>output_MAC_0_406, I407=>output_MAC_0_407, I408=>output_MAC_0_408, I409=>output_MAC_0_409, I410=>output_MAC_0_410, I411=>output_MAC_0_411, I412=>output_MAC_0_412, I413=>output_MAC_0_413, I414=>output_MAC_0_414, I415=>output_MAC_0_415, I416=>output_MAC_0_416, I417=>output_MAC_0_417, I418=>output_MAC_0_418, I419=>output_MAC_0_419, I420=>output_MAC_0_420, I421=>output_MAC_0_421, I422=>output_MAC_0_422, I423=>output_MAC_0_423, I424=>output_MAC_0_424, I425=>output_MAC_0_425, I426=>output_MAC_0_426, I427=>output_MAC_0_427, I428=>output_MAC_0_428, I429=>output_MAC_0_429, I430=>output_MAC_0_430, I431=>output_MAC_0_431, I432=>output_MAC_0_432, I433=>output_MAC_0_433, I434=>output_MAC_0_434, I435=>output_MAC_0_435, I436=>output_MAC_0_436, I437=>output_MAC_0_437, I438=>output_MAC_0_438, I439=>output_MAC_0_439, I440=>output_MAC_0_440, I441=>output_MAC_0_441, I442=>output_MAC_0_442, I443=>output_MAC_0_443, I444=>output_MAC_0_444, I445=>output_MAC_0_445, I446=>output_MAC_0_446, I447=>output_MAC_0_447, I448=>output_MAC_0_448, I449=>output_MAC_0_449, I450=>output_MAC_0_450, I451=>output_MAC_0_451, I452=>output_MAC_0_452, I453=>output_MAC_0_453, I454=>output_MAC_0_454, I455=>output_MAC_0_455, I456=>output_MAC_0_456, I457=>output_MAC_0_457, I458=>output_MAC_0_458, I459=>output_MAC_0_459, I460=>output_MAC_0_460, I461=>output_MAC_0_461, I462=>output_MAC_0_462, I463=>output_MAC_0_463, I464=>output_MAC_0_464, I465=>output_MAC_0_465, I466=>output_MAC_0_466, I467=>output_MAC_0_467, I468=>output_MAC_0_468, I469=>output_MAC_0_469, I470=>output_MAC_0_470, I471=>output_MAC_0_471, I472=>output_MAC_0_472, I473=>output_MAC_0_473, I474=>output_MAC_0_474, I475=>output_MAC_0_475, I476=>output_MAC_0_476, I477=>output_MAC_0_477, I478=>output_MAC_0_478, I479=>output_MAC_0_479, I480=>output_MAC_0_480, I481=>output_MAC_0_481, I482=>output_MAC_0_482, I483=>output_MAC_0_483, I484=>output_MAC_0_484, I485=>output_MAC_0_485, I486=>output_MAC_0_486, I487=>output_MAC_0_487, I488=>output_MAC_0_488, I489=>output_MAC_0_489, I490=>output_MAC_0_490, I491=>output_MAC_0_491, I492=>output_MAC_0_492, I493=>output_MAC_0_493, I494=>output_MAC_0_494, I495=>output_MAC_0_495, I496=>output_MAC_0_496, I497=>output_MAC_0_497, I498=>output_MAC_0_498, I499=>output_MAC_0_499, I500=>output_MAC_0_500, I501=>output_MAC_0_501, I502=>output_MAC_0_502, I503=>output_MAC_0_503, I504=>output_MAC_0_504, I505=>output_MAC_0_505, I506=>output_MAC_0_506, I507=>output_MAC_0_507, I508=>output_MAC_0_508, I509=>output_MAC_0_509, I510=>output_MAC_0_510, I511=>output_MAC_0_511, I512=>output_MAC_0_512, I513=>output_MAC_0_513, I514=>output_MAC_0_514, I515=>output_MAC_0_515, I516=>output_MAC_0_516, I517=>output_MAC_0_517, I518=>output_MAC_0_518, I519=>output_MAC_0_519, I520=>output_MAC_0_520, I521=>output_MAC_0_521, I522=>output_MAC_0_522, I523=>output_MAC_0_523, I524=>output_MAC_0_524, I525=>output_MAC_0_525, I526=>output_MAC_0_526, I527=>output_MAC_0_527, I528=>output_MAC_0_528, I529=>output_MAC_0_529, I530=>output_MAC_0_530, I531=>output_MAC_0_531, I532=>output_MAC_0_532, I533=>output_MAC_0_533, I534=>output_MAC_0_534, I535=>output_MAC_0_535, I536=>output_MAC_0_536, I537=>output_MAC_0_537, I538=>output_MAC_0_538, I539=>output_MAC_0_539, I540=>output_MAC_0_540, I541=>output_MAC_0_541, I542=>output_MAC_0_542, I543=>output_MAC_0_543, I544=>output_MAC_0_544, I545=>output_MAC_0_545, I546=>output_MAC_0_546, I547=>output_MAC_0_547, I548=>output_MAC_0_548, I549=>output_MAC_0_549, I550=>output_MAC_0_550, I551=>output_MAC_0_551, I552=>output_MAC_0_552, I553=>output_MAC_0_553, I554=>output_MAC_0_554, I555=>output_MAC_0_555, I556=>output_MAC_0_556, I557=>output_MAC_0_557, I558=>output_MAC_0_558, I559=>output_MAC_0_559, I560=>output_MAC_0_560, I561=>output_MAC_0_561, I562=>output_MAC_0_562, I563=>output_MAC_0_563, I564=>output_MAC_0_564, I565=>output_MAC_0_565, I566=>output_MAC_0_566, I567=>output_MAC_0_567, I568=>output_MAC_0_568, I569=>output_MAC_0_569, I570=>output_MAC_0_570, I571=>output_MAC_0_571, I572=>output_MAC_0_572, I573=>output_MAC_0_573, I574=>output_MAC_0_574, I575=>output_MAC_0_575, I576=>output_MAC_0_576, I577=>output_MAC_0_577, I578=>output_MAC_0_578, I579=>output_MAC_0_579, I580=>output_MAC_0_580, I581=>output_MAC_0_581, I582=>output_MAC_0_582, I583=>output_MAC_0_583, I584=>output_MAC_0_584, I585=>output_MAC_0_585, I586=>output_MAC_0_586, I587=>output_MAC_0_587, I588=>output_MAC_0_588, I589=>output_MAC_0_589, I590=>output_MAC_0_590, I591=>output_MAC_0_591, I592=>output_MAC_0_592, I593=>output_MAC_0_593, I594=>output_MAC_0_594, I595=>output_MAC_0_595, I596=>output_MAC_0_596, I597=>output_MAC_0_597, I598=>output_MAC_0_598, I599=>output_MAC_0_599, I600=>output_MAC_0_600, I601=>output_MAC_0_601, I602=>output_MAC_0_602, I603=>output_MAC_0_603, I604=>output_MAC_0_604, I605=>output_MAC_0_605, I606=>output_MAC_0_606, I607=>output_MAC_0_607, I608=>output_MAC_0_608, I609=>output_MAC_0_609, I610=>output_MAC_0_610, I611=>output_MAC_0_611, I612=>output_MAC_0_612, I613=>output_MAC_0_613, I614=>output_MAC_0_614, I615=>output_MAC_0_615, I616=>output_MAC_0_616, I617=>output_MAC_0_617, I618=>output_MAC_0_618, I619=>output_MAC_0_619, I620=>output_MAC_0_620, I621=>output_MAC_0_621, I622=>output_MAC_0_622, I623=>output_MAC_0_623, I624=>output_MAC_0_624, I625=>output_MAC_0_625, I626=>output_MAC_0_626, I627=>output_MAC_0_627, I628=>output_MAC_0_628, I629=>output_MAC_0_629, I630=>output_MAC_0_630, I631=>output_MAC_0_631, I632=>output_MAC_0_632, I633=>output_MAC_0_633, I634=>output_MAC_0_634, I635=>output_MAC_0_635, I636=>output_MAC_0_636, I637=>output_MAC_0_637, I638=>output_MAC_0_638, I639=>output_MAC_0_639, I640=>output_MAC_0_640, I641=>output_MAC_0_641, I642=>output_MAC_0_642, I643=>output_MAC_0_643, I644=>output_MAC_0_644, I645=>output_MAC_0_645, I646=>output_MAC_0_646, I647=>output_MAC_0_647, I648=>output_MAC_0_648, I649=>output_MAC_0_649, I650=>output_MAC_0_650, I651=>output_MAC_0_651, I652=>output_MAC_0_652, I653=>output_MAC_0_653, I654=>output_MAC_0_654, I655=>output_MAC_0_655, I656=>output_MAC_0_656, I657=>output_MAC_0_657, I658=>output_MAC_0_658, I659=>output_MAC_0_659, I660=>output_MAC_0_660, I661=>output_MAC_0_661, I662=>output_MAC_0_662, I663=>output_MAC_0_663, I664=>output_MAC_0_664, I665=>output_MAC_0_665, I666=>output_MAC_0_666, I667=>output_MAC_0_667, I668=>output_MAC_0_668, I669=>output_MAC_0_669, I670=>output_MAC_0_670, I671=>output_MAC_0_671, I672=>output_MAC_0_672, I673=>output_MAC_0_673, I674=>output_MAC_0_674, I675=>output_MAC_0_675, I676=>output_MAC_0_676, I677=>output_MAC_0_677, I678=>output_MAC_0_678, I679=>output_MAC_0_679, I680=>output_MAC_0_680, I681=>output_MAC_0_681, I682=>output_MAC_0_682, I683=>output_MAC_0_683, I684=>output_MAC_0_684, I685=>output_MAC_0_685, I686=>output_MAC_0_686, I687=>output_MAC_0_687, I688=>output_MAC_0_688, I689=>output_MAC_0_689, I690=>output_MAC_0_690, I691=>output_MAC_0_691, I692=>output_MAC_0_692, I693=>output_MAC_0_693, I694=>output_MAC_0_694, I695=>output_MAC_0_695, I696=>output_MAC_0_696, I697=>output_MAC_0_697, I698=>output_MAC_0_698, I699=>output_MAC_0_699, I700=>output_MAC_0_700, I701=>output_MAC_0_701, I702=>output_MAC_0_702, I703=>output_MAC_0_703, I704=>output_MAC_0_704, I705=>output_MAC_0_705, I706=>output_MAC_0_706, I707=>output_MAC_0_707, I708=>output_MAC_0_708, I709=>output_MAC_0_709, I710=>output_MAC_0_710, I711=>output_MAC_0_711, I712=>output_MAC_0_712, I713=>output_MAC_0_713, I714=>output_MAC_0_714, I715=>output_MAC_0_715, I716=>output_MAC_0_716, I717=>output_MAC_0_717, I718=>output_MAC_0_718, I719=>output_MAC_0_719, I720=>output_MAC_0_720, I721=>output_MAC_0_721, I722=>output_MAC_0_722, I723=>output_MAC_0_723, I724=>output_MAC_0_724, I725=>output_MAC_0_725, I726=>output_MAC_0_726, I727=>output_MAC_0_727, I728=>output_MAC_0_728, I729=>output_MAC_0_729, I730=>output_MAC_0_730, I731=>output_MAC_0_731, I732=>output_MAC_0_732, I733=>output_MAC_0_733, I734=>output_MAC_0_734, I735=>output_MAC_0_735, I736=>output_MAC_0_736, I737=>output_MAC_0_737, I738=>output_MAC_0_738, I739=>output_MAC_0_739, I740=>output_MAC_0_740, I741=>output_MAC_0_741, I742=>output_MAC_0_742, I743=>output_MAC_0_743, I744=>output_MAC_0_744, I745=>output_MAC_0_745, I746=>output_MAC_0_746, I747=>output_MAC_0_747, I748=>output_MAC_0_748, I749=>output_MAC_0_749, I750=>output_MAC_0_750, I751=>output_MAC_0_751, I752=>output_MAC_0_752, I753=>output_MAC_0_753, I754=>output_MAC_0_754, I755=>output_MAC_0_755, I756=>output_MAC_0_756, I757=>output_MAC_0_757, I758=>output_MAC_0_758, I759=>output_MAC_0_759, I760=>output_MAC_0_760, I761=>output_MAC_0_761, I762=>output_MAC_0_762, I763=>output_MAC_0_763, I764=>output_MAC_0_764, I765=>output_MAC_0_765, I766=>output_MAC_0_766, I767=>output_MAC_0_767, 
		SEL_mux=>SEL_mux, O=>output_row_0);

	mux_row_1: mux_768to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_1_0, I1=>output_MAC_1_1, I2=>output_MAC_1_2, I3=>output_MAC_1_3, I4=>output_MAC_1_4, I5=>output_MAC_1_5, I6=>output_MAC_1_6, I7=>output_MAC_1_7, I8=>output_MAC_1_8, I9=>output_MAC_1_9, I10=>output_MAC_1_10, I11=>output_MAC_1_11, I12=>output_MAC_1_12, I13=>output_MAC_1_13, I14=>output_MAC_1_14, I15=>output_MAC_1_15, I16=>output_MAC_1_16, I17=>output_MAC_1_17, I18=>output_MAC_1_18, I19=>output_MAC_1_19, I20=>output_MAC_1_20, I21=>output_MAC_1_21, I22=>output_MAC_1_22, I23=>output_MAC_1_23, I24=>output_MAC_1_24, I25=>output_MAC_1_25, I26=>output_MAC_1_26, I27=>output_MAC_1_27, I28=>output_MAC_1_28, I29=>output_MAC_1_29, I30=>output_MAC_1_30, I31=>output_MAC_1_31, I32=>output_MAC_1_32, I33=>output_MAC_1_33, I34=>output_MAC_1_34, I35=>output_MAC_1_35, I36=>output_MAC_1_36, I37=>output_MAC_1_37, I38=>output_MAC_1_38, I39=>output_MAC_1_39, I40=>output_MAC_1_40, I41=>output_MAC_1_41, I42=>output_MAC_1_42, I43=>output_MAC_1_43, I44=>output_MAC_1_44, I45=>output_MAC_1_45, I46=>output_MAC_1_46, I47=>output_MAC_1_47, I48=>output_MAC_1_48, I49=>output_MAC_1_49, I50=>output_MAC_1_50, I51=>output_MAC_1_51, I52=>output_MAC_1_52, I53=>output_MAC_1_53, I54=>output_MAC_1_54, I55=>output_MAC_1_55, I56=>output_MAC_1_56, I57=>output_MAC_1_57, I58=>output_MAC_1_58, I59=>output_MAC_1_59, I60=>output_MAC_1_60, I61=>output_MAC_1_61, I62=>output_MAC_1_62, I63=>output_MAC_1_63, I64=>output_MAC_1_64, I65=>output_MAC_1_65, I66=>output_MAC_1_66, I67=>output_MAC_1_67, I68=>output_MAC_1_68, I69=>output_MAC_1_69, I70=>output_MAC_1_70, I71=>output_MAC_1_71, I72=>output_MAC_1_72, I73=>output_MAC_1_73, I74=>output_MAC_1_74, I75=>output_MAC_1_75, I76=>output_MAC_1_76, I77=>output_MAC_1_77, I78=>output_MAC_1_78, I79=>output_MAC_1_79, I80=>output_MAC_1_80, I81=>output_MAC_1_81, I82=>output_MAC_1_82, I83=>output_MAC_1_83, I84=>output_MAC_1_84, I85=>output_MAC_1_85, I86=>output_MAC_1_86, I87=>output_MAC_1_87, I88=>output_MAC_1_88, I89=>output_MAC_1_89, I90=>output_MAC_1_90, I91=>output_MAC_1_91, I92=>output_MAC_1_92, I93=>output_MAC_1_93, I94=>output_MAC_1_94, I95=>output_MAC_1_95, I96=>output_MAC_1_96, I97=>output_MAC_1_97, I98=>output_MAC_1_98, I99=>output_MAC_1_99, I100=>output_MAC_1_100, I101=>output_MAC_1_101, I102=>output_MAC_1_102, I103=>output_MAC_1_103, I104=>output_MAC_1_104, I105=>output_MAC_1_105, I106=>output_MAC_1_106, I107=>output_MAC_1_107, I108=>output_MAC_1_108, I109=>output_MAC_1_109, I110=>output_MAC_1_110, I111=>output_MAC_1_111, I112=>output_MAC_1_112, I113=>output_MAC_1_113, I114=>output_MAC_1_114, I115=>output_MAC_1_115, I116=>output_MAC_1_116, I117=>output_MAC_1_117, I118=>output_MAC_1_118, I119=>output_MAC_1_119, I120=>output_MAC_1_120, I121=>output_MAC_1_121, I122=>output_MAC_1_122, I123=>output_MAC_1_123, I124=>output_MAC_1_124, I125=>output_MAC_1_125, I126=>output_MAC_1_126, I127=>output_MAC_1_127, I128=>output_MAC_1_128, I129=>output_MAC_1_129, I130=>output_MAC_1_130, I131=>output_MAC_1_131, I132=>output_MAC_1_132, I133=>output_MAC_1_133, I134=>output_MAC_1_134, I135=>output_MAC_1_135, I136=>output_MAC_1_136, I137=>output_MAC_1_137, I138=>output_MAC_1_138, I139=>output_MAC_1_139, I140=>output_MAC_1_140, I141=>output_MAC_1_141, I142=>output_MAC_1_142, I143=>output_MAC_1_143, I144=>output_MAC_1_144, I145=>output_MAC_1_145, I146=>output_MAC_1_146, I147=>output_MAC_1_147, I148=>output_MAC_1_148, I149=>output_MAC_1_149, I150=>output_MAC_1_150, I151=>output_MAC_1_151, I152=>output_MAC_1_152, I153=>output_MAC_1_153, I154=>output_MAC_1_154, I155=>output_MAC_1_155, I156=>output_MAC_1_156, I157=>output_MAC_1_157, I158=>output_MAC_1_158, I159=>output_MAC_1_159, I160=>output_MAC_1_160, I161=>output_MAC_1_161, I162=>output_MAC_1_162, I163=>output_MAC_1_163, I164=>output_MAC_1_164, I165=>output_MAC_1_165, I166=>output_MAC_1_166, I167=>output_MAC_1_167, I168=>output_MAC_1_168, I169=>output_MAC_1_169, I170=>output_MAC_1_170, I171=>output_MAC_1_171, I172=>output_MAC_1_172, I173=>output_MAC_1_173, I174=>output_MAC_1_174, I175=>output_MAC_1_175, I176=>output_MAC_1_176, I177=>output_MAC_1_177, I178=>output_MAC_1_178, I179=>output_MAC_1_179, I180=>output_MAC_1_180, I181=>output_MAC_1_181, I182=>output_MAC_1_182, I183=>output_MAC_1_183, I184=>output_MAC_1_184, I185=>output_MAC_1_185, I186=>output_MAC_1_186, I187=>output_MAC_1_187, I188=>output_MAC_1_188, I189=>output_MAC_1_189, I190=>output_MAC_1_190, I191=>output_MAC_1_191, I192=>output_MAC_1_192, I193=>output_MAC_1_193, I194=>output_MAC_1_194, I195=>output_MAC_1_195, I196=>output_MAC_1_196, I197=>output_MAC_1_197, I198=>output_MAC_1_198, I199=>output_MAC_1_199, I200=>output_MAC_1_200, I201=>output_MAC_1_201, I202=>output_MAC_1_202, I203=>output_MAC_1_203, I204=>output_MAC_1_204, I205=>output_MAC_1_205, I206=>output_MAC_1_206, I207=>output_MAC_1_207, I208=>output_MAC_1_208, I209=>output_MAC_1_209, I210=>output_MAC_1_210, I211=>output_MAC_1_211, I212=>output_MAC_1_212, I213=>output_MAC_1_213, I214=>output_MAC_1_214, I215=>output_MAC_1_215, I216=>output_MAC_1_216, I217=>output_MAC_1_217, I218=>output_MAC_1_218, I219=>output_MAC_1_219, I220=>output_MAC_1_220, I221=>output_MAC_1_221, I222=>output_MAC_1_222, I223=>output_MAC_1_223, I224=>output_MAC_1_224, I225=>output_MAC_1_225, I226=>output_MAC_1_226, I227=>output_MAC_1_227, I228=>output_MAC_1_228, I229=>output_MAC_1_229, I230=>output_MAC_1_230, I231=>output_MAC_1_231, I232=>output_MAC_1_232, I233=>output_MAC_1_233, I234=>output_MAC_1_234, I235=>output_MAC_1_235, I236=>output_MAC_1_236, I237=>output_MAC_1_237, I238=>output_MAC_1_238, I239=>output_MAC_1_239, I240=>output_MAC_1_240, I241=>output_MAC_1_241, I242=>output_MAC_1_242, I243=>output_MAC_1_243, I244=>output_MAC_1_244, I245=>output_MAC_1_245, I246=>output_MAC_1_246, I247=>output_MAC_1_247, I248=>output_MAC_1_248, I249=>output_MAC_1_249, I250=>output_MAC_1_250, I251=>output_MAC_1_251, I252=>output_MAC_1_252, I253=>output_MAC_1_253, I254=>output_MAC_1_254, I255=>output_MAC_1_255, I256=>output_MAC_1_256, I257=>output_MAC_1_257, I258=>output_MAC_1_258, I259=>output_MAC_1_259, I260=>output_MAC_1_260, I261=>output_MAC_1_261, I262=>output_MAC_1_262, I263=>output_MAC_1_263, I264=>output_MAC_1_264, I265=>output_MAC_1_265, I266=>output_MAC_1_266, I267=>output_MAC_1_267, I268=>output_MAC_1_268, I269=>output_MAC_1_269, I270=>output_MAC_1_270, I271=>output_MAC_1_271, I272=>output_MAC_1_272, I273=>output_MAC_1_273, I274=>output_MAC_1_274, I275=>output_MAC_1_275, I276=>output_MAC_1_276, I277=>output_MAC_1_277, I278=>output_MAC_1_278, I279=>output_MAC_1_279, I280=>output_MAC_1_280, I281=>output_MAC_1_281, I282=>output_MAC_1_282, I283=>output_MAC_1_283, I284=>output_MAC_1_284, I285=>output_MAC_1_285, I286=>output_MAC_1_286, I287=>output_MAC_1_287, I288=>output_MAC_1_288, I289=>output_MAC_1_289, I290=>output_MAC_1_290, I291=>output_MAC_1_291, I292=>output_MAC_1_292, I293=>output_MAC_1_293, I294=>output_MAC_1_294, I295=>output_MAC_1_295, I296=>output_MAC_1_296, I297=>output_MAC_1_297, I298=>output_MAC_1_298, I299=>output_MAC_1_299, I300=>output_MAC_1_300, I301=>output_MAC_1_301, I302=>output_MAC_1_302, I303=>output_MAC_1_303, I304=>output_MAC_1_304, I305=>output_MAC_1_305, I306=>output_MAC_1_306, I307=>output_MAC_1_307, I308=>output_MAC_1_308, I309=>output_MAC_1_309, I310=>output_MAC_1_310, I311=>output_MAC_1_311, I312=>output_MAC_1_312, I313=>output_MAC_1_313, I314=>output_MAC_1_314, I315=>output_MAC_1_315, I316=>output_MAC_1_316, I317=>output_MAC_1_317, I318=>output_MAC_1_318, I319=>output_MAC_1_319, I320=>output_MAC_1_320, I321=>output_MAC_1_321, I322=>output_MAC_1_322, I323=>output_MAC_1_323, I324=>output_MAC_1_324, I325=>output_MAC_1_325, I326=>output_MAC_1_326, I327=>output_MAC_1_327, I328=>output_MAC_1_328, I329=>output_MAC_1_329, I330=>output_MAC_1_330, I331=>output_MAC_1_331, I332=>output_MAC_1_332, I333=>output_MAC_1_333, I334=>output_MAC_1_334, I335=>output_MAC_1_335, I336=>output_MAC_1_336, I337=>output_MAC_1_337, I338=>output_MAC_1_338, I339=>output_MAC_1_339, I340=>output_MAC_1_340, I341=>output_MAC_1_341, I342=>output_MAC_1_342, I343=>output_MAC_1_343, I344=>output_MAC_1_344, I345=>output_MAC_1_345, I346=>output_MAC_1_346, I347=>output_MAC_1_347, I348=>output_MAC_1_348, I349=>output_MAC_1_349, I350=>output_MAC_1_350, I351=>output_MAC_1_351, I352=>output_MAC_1_352, I353=>output_MAC_1_353, I354=>output_MAC_1_354, I355=>output_MAC_1_355, I356=>output_MAC_1_356, I357=>output_MAC_1_357, I358=>output_MAC_1_358, I359=>output_MAC_1_359, I360=>output_MAC_1_360, I361=>output_MAC_1_361, I362=>output_MAC_1_362, I363=>output_MAC_1_363, I364=>output_MAC_1_364, I365=>output_MAC_1_365, I366=>output_MAC_1_366, I367=>output_MAC_1_367, I368=>output_MAC_1_368, I369=>output_MAC_1_369, I370=>output_MAC_1_370, I371=>output_MAC_1_371, I372=>output_MAC_1_372, I373=>output_MAC_1_373, I374=>output_MAC_1_374, I375=>output_MAC_1_375, I376=>output_MAC_1_376, I377=>output_MAC_1_377, I378=>output_MAC_1_378, I379=>output_MAC_1_379, I380=>output_MAC_1_380, I381=>output_MAC_1_381, I382=>output_MAC_1_382, I383=>output_MAC_1_383, I384=>output_MAC_1_384, I385=>output_MAC_1_385, I386=>output_MAC_1_386, I387=>output_MAC_1_387, I388=>output_MAC_1_388, I389=>output_MAC_1_389, I390=>output_MAC_1_390, I391=>output_MAC_1_391, I392=>output_MAC_1_392, I393=>output_MAC_1_393, I394=>output_MAC_1_394, I395=>output_MAC_1_395, I396=>output_MAC_1_396, I397=>output_MAC_1_397, I398=>output_MAC_1_398, I399=>output_MAC_1_399, I400=>output_MAC_1_400, I401=>output_MAC_1_401, I402=>output_MAC_1_402, I403=>output_MAC_1_403, I404=>output_MAC_1_404, I405=>output_MAC_1_405, I406=>output_MAC_1_406, I407=>output_MAC_1_407, I408=>output_MAC_1_408, I409=>output_MAC_1_409, I410=>output_MAC_1_410, I411=>output_MAC_1_411, I412=>output_MAC_1_412, I413=>output_MAC_1_413, I414=>output_MAC_1_414, I415=>output_MAC_1_415, I416=>output_MAC_1_416, I417=>output_MAC_1_417, I418=>output_MAC_1_418, I419=>output_MAC_1_419, I420=>output_MAC_1_420, I421=>output_MAC_1_421, I422=>output_MAC_1_422, I423=>output_MAC_1_423, I424=>output_MAC_1_424, I425=>output_MAC_1_425, I426=>output_MAC_1_426, I427=>output_MAC_1_427, I428=>output_MAC_1_428, I429=>output_MAC_1_429, I430=>output_MAC_1_430, I431=>output_MAC_1_431, I432=>output_MAC_1_432, I433=>output_MAC_1_433, I434=>output_MAC_1_434, I435=>output_MAC_1_435, I436=>output_MAC_1_436, I437=>output_MAC_1_437, I438=>output_MAC_1_438, I439=>output_MAC_1_439, I440=>output_MAC_1_440, I441=>output_MAC_1_441, I442=>output_MAC_1_442, I443=>output_MAC_1_443, I444=>output_MAC_1_444, I445=>output_MAC_1_445, I446=>output_MAC_1_446, I447=>output_MAC_1_447, I448=>output_MAC_1_448, I449=>output_MAC_1_449, I450=>output_MAC_1_450, I451=>output_MAC_1_451, I452=>output_MAC_1_452, I453=>output_MAC_1_453, I454=>output_MAC_1_454, I455=>output_MAC_1_455, I456=>output_MAC_1_456, I457=>output_MAC_1_457, I458=>output_MAC_1_458, I459=>output_MAC_1_459, I460=>output_MAC_1_460, I461=>output_MAC_1_461, I462=>output_MAC_1_462, I463=>output_MAC_1_463, I464=>output_MAC_1_464, I465=>output_MAC_1_465, I466=>output_MAC_1_466, I467=>output_MAC_1_467, I468=>output_MAC_1_468, I469=>output_MAC_1_469, I470=>output_MAC_1_470, I471=>output_MAC_1_471, I472=>output_MAC_1_472, I473=>output_MAC_1_473, I474=>output_MAC_1_474, I475=>output_MAC_1_475, I476=>output_MAC_1_476, I477=>output_MAC_1_477, I478=>output_MAC_1_478, I479=>output_MAC_1_479, I480=>output_MAC_1_480, I481=>output_MAC_1_481, I482=>output_MAC_1_482, I483=>output_MAC_1_483, I484=>output_MAC_1_484, I485=>output_MAC_1_485, I486=>output_MAC_1_486, I487=>output_MAC_1_487, I488=>output_MAC_1_488, I489=>output_MAC_1_489, I490=>output_MAC_1_490, I491=>output_MAC_1_491, I492=>output_MAC_1_492, I493=>output_MAC_1_493, I494=>output_MAC_1_494, I495=>output_MAC_1_495, I496=>output_MAC_1_496, I497=>output_MAC_1_497, I498=>output_MAC_1_498, I499=>output_MAC_1_499, I500=>output_MAC_1_500, I501=>output_MAC_1_501, I502=>output_MAC_1_502, I503=>output_MAC_1_503, I504=>output_MAC_1_504, I505=>output_MAC_1_505, I506=>output_MAC_1_506, I507=>output_MAC_1_507, I508=>output_MAC_1_508, I509=>output_MAC_1_509, I510=>output_MAC_1_510, I511=>output_MAC_1_511, I512=>output_MAC_1_512, I513=>output_MAC_1_513, I514=>output_MAC_1_514, I515=>output_MAC_1_515, I516=>output_MAC_1_516, I517=>output_MAC_1_517, I518=>output_MAC_1_518, I519=>output_MAC_1_519, I520=>output_MAC_1_520, I521=>output_MAC_1_521, I522=>output_MAC_1_522, I523=>output_MAC_1_523, I524=>output_MAC_1_524, I525=>output_MAC_1_525, I526=>output_MAC_1_526, I527=>output_MAC_1_527, I528=>output_MAC_1_528, I529=>output_MAC_1_529, I530=>output_MAC_1_530, I531=>output_MAC_1_531, I532=>output_MAC_1_532, I533=>output_MAC_1_533, I534=>output_MAC_1_534, I535=>output_MAC_1_535, I536=>output_MAC_1_536, I537=>output_MAC_1_537, I538=>output_MAC_1_538, I539=>output_MAC_1_539, I540=>output_MAC_1_540, I541=>output_MAC_1_541, I542=>output_MAC_1_542, I543=>output_MAC_1_543, I544=>output_MAC_1_544, I545=>output_MAC_1_545, I546=>output_MAC_1_546, I547=>output_MAC_1_547, I548=>output_MAC_1_548, I549=>output_MAC_1_549, I550=>output_MAC_1_550, I551=>output_MAC_1_551, I552=>output_MAC_1_552, I553=>output_MAC_1_553, I554=>output_MAC_1_554, I555=>output_MAC_1_555, I556=>output_MAC_1_556, I557=>output_MAC_1_557, I558=>output_MAC_1_558, I559=>output_MAC_1_559, I560=>output_MAC_1_560, I561=>output_MAC_1_561, I562=>output_MAC_1_562, I563=>output_MAC_1_563, I564=>output_MAC_1_564, I565=>output_MAC_1_565, I566=>output_MAC_1_566, I567=>output_MAC_1_567, I568=>output_MAC_1_568, I569=>output_MAC_1_569, I570=>output_MAC_1_570, I571=>output_MAC_1_571, I572=>output_MAC_1_572, I573=>output_MAC_1_573, I574=>output_MAC_1_574, I575=>output_MAC_1_575, I576=>output_MAC_1_576, I577=>output_MAC_1_577, I578=>output_MAC_1_578, I579=>output_MAC_1_579, I580=>output_MAC_1_580, I581=>output_MAC_1_581, I582=>output_MAC_1_582, I583=>output_MAC_1_583, I584=>output_MAC_1_584, I585=>output_MAC_1_585, I586=>output_MAC_1_586, I587=>output_MAC_1_587, I588=>output_MAC_1_588, I589=>output_MAC_1_589, I590=>output_MAC_1_590, I591=>output_MAC_1_591, I592=>output_MAC_1_592, I593=>output_MAC_1_593, I594=>output_MAC_1_594, I595=>output_MAC_1_595, I596=>output_MAC_1_596, I597=>output_MAC_1_597, I598=>output_MAC_1_598, I599=>output_MAC_1_599, I600=>output_MAC_1_600, I601=>output_MAC_1_601, I602=>output_MAC_1_602, I603=>output_MAC_1_603, I604=>output_MAC_1_604, I605=>output_MAC_1_605, I606=>output_MAC_1_606, I607=>output_MAC_1_607, I608=>output_MAC_1_608, I609=>output_MAC_1_609, I610=>output_MAC_1_610, I611=>output_MAC_1_611, I612=>output_MAC_1_612, I613=>output_MAC_1_613, I614=>output_MAC_1_614, I615=>output_MAC_1_615, I616=>output_MAC_1_616, I617=>output_MAC_1_617, I618=>output_MAC_1_618, I619=>output_MAC_1_619, I620=>output_MAC_1_620, I621=>output_MAC_1_621, I622=>output_MAC_1_622, I623=>output_MAC_1_623, I624=>output_MAC_1_624, I625=>output_MAC_1_625, I626=>output_MAC_1_626, I627=>output_MAC_1_627, I628=>output_MAC_1_628, I629=>output_MAC_1_629, I630=>output_MAC_1_630, I631=>output_MAC_1_631, I632=>output_MAC_1_632, I633=>output_MAC_1_633, I634=>output_MAC_1_634, I635=>output_MAC_1_635, I636=>output_MAC_1_636, I637=>output_MAC_1_637, I638=>output_MAC_1_638, I639=>output_MAC_1_639, I640=>output_MAC_1_640, I641=>output_MAC_1_641, I642=>output_MAC_1_642, I643=>output_MAC_1_643, I644=>output_MAC_1_644, I645=>output_MAC_1_645, I646=>output_MAC_1_646, I647=>output_MAC_1_647, I648=>output_MAC_1_648, I649=>output_MAC_1_649, I650=>output_MAC_1_650, I651=>output_MAC_1_651, I652=>output_MAC_1_652, I653=>output_MAC_1_653, I654=>output_MAC_1_654, I655=>output_MAC_1_655, I656=>output_MAC_1_656, I657=>output_MAC_1_657, I658=>output_MAC_1_658, I659=>output_MAC_1_659, I660=>output_MAC_1_660, I661=>output_MAC_1_661, I662=>output_MAC_1_662, I663=>output_MAC_1_663, I664=>output_MAC_1_664, I665=>output_MAC_1_665, I666=>output_MAC_1_666, I667=>output_MAC_1_667, I668=>output_MAC_1_668, I669=>output_MAC_1_669, I670=>output_MAC_1_670, I671=>output_MAC_1_671, I672=>output_MAC_1_672, I673=>output_MAC_1_673, I674=>output_MAC_1_674, I675=>output_MAC_1_675, I676=>output_MAC_1_676, I677=>output_MAC_1_677, I678=>output_MAC_1_678, I679=>output_MAC_1_679, I680=>output_MAC_1_680, I681=>output_MAC_1_681, I682=>output_MAC_1_682, I683=>output_MAC_1_683, I684=>output_MAC_1_684, I685=>output_MAC_1_685, I686=>output_MAC_1_686, I687=>output_MAC_1_687, I688=>output_MAC_1_688, I689=>output_MAC_1_689, I690=>output_MAC_1_690, I691=>output_MAC_1_691, I692=>output_MAC_1_692, I693=>output_MAC_1_693, I694=>output_MAC_1_694, I695=>output_MAC_1_695, I696=>output_MAC_1_696, I697=>output_MAC_1_697, I698=>output_MAC_1_698, I699=>output_MAC_1_699, I700=>output_MAC_1_700, I701=>output_MAC_1_701, I702=>output_MAC_1_702, I703=>output_MAC_1_703, I704=>output_MAC_1_704, I705=>output_MAC_1_705, I706=>output_MAC_1_706, I707=>output_MAC_1_707, I708=>output_MAC_1_708, I709=>output_MAC_1_709, I710=>output_MAC_1_710, I711=>output_MAC_1_711, I712=>output_MAC_1_712, I713=>output_MAC_1_713, I714=>output_MAC_1_714, I715=>output_MAC_1_715, I716=>output_MAC_1_716, I717=>output_MAC_1_717, I718=>output_MAC_1_718, I719=>output_MAC_1_719, I720=>output_MAC_1_720, I721=>output_MAC_1_721, I722=>output_MAC_1_722, I723=>output_MAC_1_723, I724=>output_MAC_1_724, I725=>output_MAC_1_725, I726=>output_MAC_1_726, I727=>output_MAC_1_727, I728=>output_MAC_1_728, I729=>output_MAC_1_729, I730=>output_MAC_1_730, I731=>output_MAC_1_731, I732=>output_MAC_1_732, I733=>output_MAC_1_733, I734=>output_MAC_1_734, I735=>output_MAC_1_735, I736=>output_MAC_1_736, I737=>output_MAC_1_737, I738=>output_MAC_1_738, I739=>output_MAC_1_739, I740=>output_MAC_1_740, I741=>output_MAC_1_741, I742=>output_MAC_1_742, I743=>output_MAC_1_743, I744=>output_MAC_1_744, I745=>output_MAC_1_745, I746=>output_MAC_1_746, I747=>output_MAC_1_747, I748=>output_MAC_1_748, I749=>output_MAC_1_749, I750=>output_MAC_1_750, I751=>output_MAC_1_751, I752=>output_MAC_1_752, I753=>output_MAC_1_753, I754=>output_MAC_1_754, I755=>output_MAC_1_755, I756=>output_MAC_1_756, I757=>output_MAC_1_757, I758=>output_MAC_1_758, I759=>output_MAC_1_759, I760=>output_MAC_1_760, I761=>output_MAC_1_761, I762=>output_MAC_1_762, I763=>output_MAC_1_763, I764=>output_MAC_1_764, I765=>output_MAC_1_765, I766=>output_MAC_1_766, I767=>output_MAC_1_767, 
		SEL_mux=>SEL_mux, O=>output_row_1);

	mux_row_2: mux_768to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_2_0, I1=>output_MAC_2_1, I2=>output_MAC_2_2, I3=>output_MAC_2_3, I4=>output_MAC_2_4, I5=>output_MAC_2_5, I6=>output_MAC_2_6, I7=>output_MAC_2_7, I8=>output_MAC_2_8, I9=>output_MAC_2_9, I10=>output_MAC_2_10, I11=>output_MAC_2_11, I12=>output_MAC_2_12, I13=>output_MAC_2_13, I14=>output_MAC_2_14, I15=>output_MAC_2_15, I16=>output_MAC_2_16, I17=>output_MAC_2_17, I18=>output_MAC_2_18, I19=>output_MAC_2_19, I20=>output_MAC_2_20, I21=>output_MAC_2_21, I22=>output_MAC_2_22, I23=>output_MAC_2_23, I24=>output_MAC_2_24, I25=>output_MAC_2_25, I26=>output_MAC_2_26, I27=>output_MAC_2_27, I28=>output_MAC_2_28, I29=>output_MAC_2_29, I30=>output_MAC_2_30, I31=>output_MAC_2_31, I32=>output_MAC_2_32, I33=>output_MAC_2_33, I34=>output_MAC_2_34, I35=>output_MAC_2_35, I36=>output_MAC_2_36, I37=>output_MAC_2_37, I38=>output_MAC_2_38, I39=>output_MAC_2_39, I40=>output_MAC_2_40, I41=>output_MAC_2_41, I42=>output_MAC_2_42, I43=>output_MAC_2_43, I44=>output_MAC_2_44, I45=>output_MAC_2_45, I46=>output_MAC_2_46, I47=>output_MAC_2_47, I48=>output_MAC_2_48, I49=>output_MAC_2_49, I50=>output_MAC_2_50, I51=>output_MAC_2_51, I52=>output_MAC_2_52, I53=>output_MAC_2_53, I54=>output_MAC_2_54, I55=>output_MAC_2_55, I56=>output_MAC_2_56, I57=>output_MAC_2_57, I58=>output_MAC_2_58, I59=>output_MAC_2_59, I60=>output_MAC_2_60, I61=>output_MAC_2_61, I62=>output_MAC_2_62, I63=>output_MAC_2_63, I64=>output_MAC_2_64, I65=>output_MAC_2_65, I66=>output_MAC_2_66, I67=>output_MAC_2_67, I68=>output_MAC_2_68, I69=>output_MAC_2_69, I70=>output_MAC_2_70, I71=>output_MAC_2_71, I72=>output_MAC_2_72, I73=>output_MAC_2_73, I74=>output_MAC_2_74, I75=>output_MAC_2_75, I76=>output_MAC_2_76, I77=>output_MAC_2_77, I78=>output_MAC_2_78, I79=>output_MAC_2_79, I80=>output_MAC_2_80, I81=>output_MAC_2_81, I82=>output_MAC_2_82, I83=>output_MAC_2_83, I84=>output_MAC_2_84, I85=>output_MAC_2_85, I86=>output_MAC_2_86, I87=>output_MAC_2_87, I88=>output_MAC_2_88, I89=>output_MAC_2_89, I90=>output_MAC_2_90, I91=>output_MAC_2_91, I92=>output_MAC_2_92, I93=>output_MAC_2_93, I94=>output_MAC_2_94, I95=>output_MAC_2_95, I96=>output_MAC_2_96, I97=>output_MAC_2_97, I98=>output_MAC_2_98, I99=>output_MAC_2_99, I100=>output_MAC_2_100, I101=>output_MAC_2_101, I102=>output_MAC_2_102, I103=>output_MAC_2_103, I104=>output_MAC_2_104, I105=>output_MAC_2_105, I106=>output_MAC_2_106, I107=>output_MAC_2_107, I108=>output_MAC_2_108, I109=>output_MAC_2_109, I110=>output_MAC_2_110, I111=>output_MAC_2_111, I112=>output_MAC_2_112, I113=>output_MAC_2_113, I114=>output_MAC_2_114, I115=>output_MAC_2_115, I116=>output_MAC_2_116, I117=>output_MAC_2_117, I118=>output_MAC_2_118, I119=>output_MAC_2_119, I120=>output_MAC_2_120, I121=>output_MAC_2_121, I122=>output_MAC_2_122, I123=>output_MAC_2_123, I124=>output_MAC_2_124, I125=>output_MAC_2_125, I126=>output_MAC_2_126, I127=>output_MAC_2_127, I128=>output_MAC_2_128, I129=>output_MAC_2_129, I130=>output_MAC_2_130, I131=>output_MAC_2_131, I132=>output_MAC_2_132, I133=>output_MAC_2_133, I134=>output_MAC_2_134, I135=>output_MAC_2_135, I136=>output_MAC_2_136, I137=>output_MAC_2_137, I138=>output_MAC_2_138, I139=>output_MAC_2_139, I140=>output_MAC_2_140, I141=>output_MAC_2_141, I142=>output_MAC_2_142, I143=>output_MAC_2_143, I144=>output_MAC_2_144, I145=>output_MAC_2_145, I146=>output_MAC_2_146, I147=>output_MAC_2_147, I148=>output_MAC_2_148, I149=>output_MAC_2_149, I150=>output_MAC_2_150, I151=>output_MAC_2_151, I152=>output_MAC_2_152, I153=>output_MAC_2_153, I154=>output_MAC_2_154, I155=>output_MAC_2_155, I156=>output_MAC_2_156, I157=>output_MAC_2_157, I158=>output_MAC_2_158, I159=>output_MAC_2_159, I160=>output_MAC_2_160, I161=>output_MAC_2_161, I162=>output_MAC_2_162, I163=>output_MAC_2_163, I164=>output_MAC_2_164, I165=>output_MAC_2_165, I166=>output_MAC_2_166, I167=>output_MAC_2_167, I168=>output_MAC_2_168, I169=>output_MAC_2_169, I170=>output_MAC_2_170, I171=>output_MAC_2_171, I172=>output_MAC_2_172, I173=>output_MAC_2_173, I174=>output_MAC_2_174, I175=>output_MAC_2_175, I176=>output_MAC_2_176, I177=>output_MAC_2_177, I178=>output_MAC_2_178, I179=>output_MAC_2_179, I180=>output_MAC_2_180, I181=>output_MAC_2_181, I182=>output_MAC_2_182, I183=>output_MAC_2_183, I184=>output_MAC_2_184, I185=>output_MAC_2_185, I186=>output_MAC_2_186, I187=>output_MAC_2_187, I188=>output_MAC_2_188, I189=>output_MAC_2_189, I190=>output_MAC_2_190, I191=>output_MAC_2_191, I192=>output_MAC_2_192, I193=>output_MAC_2_193, I194=>output_MAC_2_194, I195=>output_MAC_2_195, I196=>output_MAC_2_196, I197=>output_MAC_2_197, I198=>output_MAC_2_198, I199=>output_MAC_2_199, I200=>output_MAC_2_200, I201=>output_MAC_2_201, I202=>output_MAC_2_202, I203=>output_MAC_2_203, I204=>output_MAC_2_204, I205=>output_MAC_2_205, I206=>output_MAC_2_206, I207=>output_MAC_2_207, I208=>output_MAC_2_208, I209=>output_MAC_2_209, I210=>output_MAC_2_210, I211=>output_MAC_2_211, I212=>output_MAC_2_212, I213=>output_MAC_2_213, I214=>output_MAC_2_214, I215=>output_MAC_2_215, I216=>output_MAC_2_216, I217=>output_MAC_2_217, I218=>output_MAC_2_218, I219=>output_MAC_2_219, I220=>output_MAC_2_220, I221=>output_MAC_2_221, I222=>output_MAC_2_222, I223=>output_MAC_2_223, I224=>output_MAC_2_224, I225=>output_MAC_2_225, I226=>output_MAC_2_226, I227=>output_MAC_2_227, I228=>output_MAC_2_228, I229=>output_MAC_2_229, I230=>output_MAC_2_230, I231=>output_MAC_2_231, I232=>output_MAC_2_232, I233=>output_MAC_2_233, I234=>output_MAC_2_234, I235=>output_MAC_2_235, I236=>output_MAC_2_236, I237=>output_MAC_2_237, I238=>output_MAC_2_238, I239=>output_MAC_2_239, I240=>output_MAC_2_240, I241=>output_MAC_2_241, I242=>output_MAC_2_242, I243=>output_MAC_2_243, I244=>output_MAC_2_244, I245=>output_MAC_2_245, I246=>output_MAC_2_246, I247=>output_MAC_2_247, I248=>output_MAC_2_248, I249=>output_MAC_2_249, I250=>output_MAC_2_250, I251=>output_MAC_2_251, I252=>output_MAC_2_252, I253=>output_MAC_2_253, I254=>output_MAC_2_254, I255=>output_MAC_2_255, I256=>output_MAC_2_256, I257=>output_MAC_2_257, I258=>output_MAC_2_258, I259=>output_MAC_2_259, I260=>output_MAC_2_260, I261=>output_MAC_2_261, I262=>output_MAC_2_262, I263=>output_MAC_2_263, I264=>output_MAC_2_264, I265=>output_MAC_2_265, I266=>output_MAC_2_266, I267=>output_MAC_2_267, I268=>output_MAC_2_268, I269=>output_MAC_2_269, I270=>output_MAC_2_270, I271=>output_MAC_2_271, I272=>output_MAC_2_272, I273=>output_MAC_2_273, I274=>output_MAC_2_274, I275=>output_MAC_2_275, I276=>output_MAC_2_276, I277=>output_MAC_2_277, I278=>output_MAC_2_278, I279=>output_MAC_2_279, I280=>output_MAC_2_280, I281=>output_MAC_2_281, I282=>output_MAC_2_282, I283=>output_MAC_2_283, I284=>output_MAC_2_284, I285=>output_MAC_2_285, I286=>output_MAC_2_286, I287=>output_MAC_2_287, I288=>output_MAC_2_288, I289=>output_MAC_2_289, I290=>output_MAC_2_290, I291=>output_MAC_2_291, I292=>output_MAC_2_292, I293=>output_MAC_2_293, I294=>output_MAC_2_294, I295=>output_MAC_2_295, I296=>output_MAC_2_296, I297=>output_MAC_2_297, I298=>output_MAC_2_298, I299=>output_MAC_2_299, I300=>output_MAC_2_300, I301=>output_MAC_2_301, I302=>output_MAC_2_302, I303=>output_MAC_2_303, I304=>output_MAC_2_304, I305=>output_MAC_2_305, I306=>output_MAC_2_306, I307=>output_MAC_2_307, I308=>output_MAC_2_308, I309=>output_MAC_2_309, I310=>output_MAC_2_310, I311=>output_MAC_2_311, I312=>output_MAC_2_312, I313=>output_MAC_2_313, I314=>output_MAC_2_314, I315=>output_MAC_2_315, I316=>output_MAC_2_316, I317=>output_MAC_2_317, I318=>output_MAC_2_318, I319=>output_MAC_2_319, I320=>output_MAC_2_320, I321=>output_MAC_2_321, I322=>output_MAC_2_322, I323=>output_MAC_2_323, I324=>output_MAC_2_324, I325=>output_MAC_2_325, I326=>output_MAC_2_326, I327=>output_MAC_2_327, I328=>output_MAC_2_328, I329=>output_MAC_2_329, I330=>output_MAC_2_330, I331=>output_MAC_2_331, I332=>output_MAC_2_332, I333=>output_MAC_2_333, I334=>output_MAC_2_334, I335=>output_MAC_2_335, I336=>output_MAC_2_336, I337=>output_MAC_2_337, I338=>output_MAC_2_338, I339=>output_MAC_2_339, I340=>output_MAC_2_340, I341=>output_MAC_2_341, I342=>output_MAC_2_342, I343=>output_MAC_2_343, I344=>output_MAC_2_344, I345=>output_MAC_2_345, I346=>output_MAC_2_346, I347=>output_MAC_2_347, I348=>output_MAC_2_348, I349=>output_MAC_2_349, I350=>output_MAC_2_350, I351=>output_MAC_2_351, I352=>output_MAC_2_352, I353=>output_MAC_2_353, I354=>output_MAC_2_354, I355=>output_MAC_2_355, I356=>output_MAC_2_356, I357=>output_MAC_2_357, I358=>output_MAC_2_358, I359=>output_MAC_2_359, I360=>output_MAC_2_360, I361=>output_MAC_2_361, I362=>output_MAC_2_362, I363=>output_MAC_2_363, I364=>output_MAC_2_364, I365=>output_MAC_2_365, I366=>output_MAC_2_366, I367=>output_MAC_2_367, I368=>output_MAC_2_368, I369=>output_MAC_2_369, I370=>output_MAC_2_370, I371=>output_MAC_2_371, I372=>output_MAC_2_372, I373=>output_MAC_2_373, I374=>output_MAC_2_374, I375=>output_MAC_2_375, I376=>output_MAC_2_376, I377=>output_MAC_2_377, I378=>output_MAC_2_378, I379=>output_MAC_2_379, I380=>output_MAC_2_380, I381=>output_MAC_2_381, I382=>output_MAC_2_382, I383=>output_MAC_2_383, I384=>output_MAC_2_384, I385=>output_MAC_2_385, I386=>output_MAC_2_386, I387=>output_MAC_2_387, I388=>output_MAC_2_388, I389=>output_MAC_2_389, I390=>output_MAC_2_390, I391=>output_MAC_2_391, I392=>output_MAC_2_392, I393=>output_MAC_2_393, I394=>output_MAC_2_394, I395=>output_MAC_2_395, I396=>output_MAC_2_396, I397=>output_MAC_2_397, I398=>output_MAC_2_398, I399=>output_MAC_2_399, I400=>output_MAC_2_400, I401=>output_MAC_2_401, I402=>output_MAC_2_402, I403=>output_MAC_2_403, I404=>output_MAC_2_404, I405=>output_MAC_2_405, I406=>output_MAC_2_406, I407=>output_MAC_2_407, I408=>output_MAC_2_408, I409=>output_MAC_2_409, I410=>output_MAC_2_410, I411=>output_MAC_2_411, I412=>output_MAC_2_412, I413=>output_MAC_2_413, I414=>output_MAC_2_414, I415=>output_MAC_2_415, I416=>output_MAC_2_416, I417=>output_MAC_2_417, I418=>output_MAC_2_418, I419=>output_MAC_2_419, I420=>output_MAC_2_420, I421=>output_MAC_2_421, I422=>output_MAC_2_422, I423=>output_MAC_2_423, I424=>output_MAC_2_424, I425=>output_MAC_2_425, I426=>output_MAC_2_426, I427=>output_MAC_2_427, I428=>output_MAC_2_428, I429=>output_MAC_2_429, I430=>output_MAC_2_430, I431=>output_MAC_2_431, I432=>output_MAC_2_432, I433=>output_MAC_2_433, I434=>output_MAC_2_434, I435=>output_MAC_2_435, I436=>output_MAC_2_436, I437=>output_MAC_2_437, I438=>output_MAC_2_438, I439=>output_MAC_2_439, I440=>output_MAC_2_440, I441=>output_MAC_2_441, I442=>output_MAC_2_442, I443=>output_MAC_2_443, I444=>output_MAC_2_444, I445=>output_MAC_2_445, I446=>output_MAC_2_446, I447=>output_MAC_2_447, I448=>output_MAC_2_448, I449=>output_MAC_2_449, I450=>output_MAC_2_450, I451=>output_MAC_2_451, I452=>output_MAC_2_452, I453=>output_MAC_2_453, I454=>output_MAC_2_454, I455=>output_MAC_2_455, I456=>output_MAC_2_456, I457=>output_MAC_2_457, I458=>output_MAC_2_458, I459=>output_MAC_2_459, I460=>output_MAC_2_460, I461=>output_MAC_2_461, I462=>output_MAC_2_462, I463=>output_MAC_2_463, I464=>output_MAC_2_464, I465=>output_MAC_2_465, I466=>output_MAC_2_466, I467=>output_MAC_2_467, I468=>output_MAC_2_468, I469=>output_MAC_2_469, I470=>output_MAC_2_470, I471=>output_MAC_2_471, I472=>output_MAC_2_472, I473=>output_MAC_2_473, I474=>output_MAC_2_474, I475=>output_MAC_2_475, I476=>output_MAC_2_476, I477=>output_MAC_2_477, I478=>output_MAC_2_478, I479=>output_MAC_2_479, I480=>output_MAC_2_480, I481=>output_MAC_2_481, I482=>output_MAC_2_482, I483=>output_MAC_2_483, I484=>output_MAC_2_484, I485=>output_MAC_2_485, I486=>output_MAC_2_486, I487=>output_MAC_2_487, I488=>output_MAC_2_488, I489=>output_MAC_2_489, I490=>output_MAC_2_490, I491=>output_MAC_2_491, I492=>output_MAC_2_492, I493=>output_MAC_2_493, I494=>output_MAC_2_494, I495=>output_MAC_2_495, I496=>output_MAC_2_496, I497=>output_MAC_2_497, I498=>output_MAC_2_498, I499=>output_MAC_2_499, I500=>output_MAC_2_500, I501=>output_MAC_2_501, I502=>output_MAC_2_502, I503=>output_MAC_2_503, I504=>output_MAC_2_504, I505=>output_MAC_2_505, I506=>output_MAC_2_506, I507=>output_MAC_2_507, I508=>output_MAC_2_508, I509=>output_MAC_2_509, I510=>output_MAC_2_510, I511=>output_MAC_2_511, I512=>output_MAC_2_512, I513=>output_MAC_2_513, I514=>output_MAC_2_514, I515=>output_MAC_2_515, I516=>output_MAC_2_516, I517=>output_MAC_2_517, I518=>output_MAC_2_518, I519=>output_MAC_2_519, I520=>output_MAC_2_520, I521=>output_MAC_2_521, I522=>output_MAC_2_522, I523=>output_MAC_2_523, I524=>output_MAC_2_524, I525=>output_MAC_2_525, I526=>output_MAC_2_526, I527=>output_MAC_2_527, I528=>output_MAC_2_528, I529=>output_MAC_2_529, I530=>output_MAC_2_530, I531=>output_MAC_2_531, I532=>output_MAC_2_532, I533=>output_MAC_2_533, I534=>output_MAC_2_534, I535=>output_MAC_2_535, I536=>output_MAC_2_536, I537=>output_MAC_2_537, I538=>output_MAC_2_538, I539=>output_MAC_2_539, I540=>output_MAC_2_540, I541=>output_MAC_2_541, I542=>output_MAC_2_542, I543=>output_MAC_2_543, I544=>output_MAC_2_544, I545=>output_MAC_2_545, I546=>output_MAC_2_546, I547=>output_MAC_2_547, I548=>output_MAC_2_548, I549=>output_MAC_2_549, I550=>output_MAC_2_550, I551=>output_MAC_2_551, I552=>output_MAC_2_552, I553=>output_MAC_2_553, I554=>output_MAC_2_554, I555=>output_MAC_2_555, I556=>output_MAC_2_556, I557=>output_MAC_2_557, I558=>output_MAC_2_558, I559=>output_MAC_2_559, I560=>output_MAC_2_560, I561=>output_MAC_2_561, I562=>output_MAC_2_562, I563=>output_MAC_2_563, I564=>output_MAC_2_564, I565=>output_MAC_2_565, I566=>output_MAC_2_566, I567=>output_MAC_2_567, I568=>output_MAC_2_568, I569=>output_MAC_2_569, I570=>output_MAC_2_570, I571=>output_MAC_2_571, I572=>output_MAC_2_572, I573=>output_MAC_2_573, I574=>output_MAC_2_574, I575=>output_MAC_2_575, I576=>output_MAC_2_576, I577=>output_MAC_2_577, I578=>output_MAC_2_578, I579=>output_MAC_2_579, I580=>output_MAC_2_580, I581=>output_MAC_2_581, I582=>output_MAC_2_582, I583=>output_MAC_2_583, I584=>output_MAC_2_584, I585=>output_MAC_2_585, I586=>output_MAC_2_586, I587=>output_MAC_2_587, I588=>output_MAC_2_588, I589=>output_MAC_2_589, I590=>output_MAC_2_590, I591=>output_MAC_2_591, I592=>output_MAC_2_592, I593=>output_MAC_2_593, I594=>output_MAC_2_594, I595=>output_MAC_2_595, I596=>output_MAC_2_596, I597=>output_MAC_2_597, I598=>output_MAC_2_598, I599=>output_MAC_2_599, I600=>output_MAC_2_600, I601=>output_MAC_2_601, I602=>output_MAC_2_602, I603=>output_MAC_2_603, I604=>output_MAC_2_604, I605=>output_MAC_2_605, I606=>output_MAC_2_606, I607=>output_MAC_2_607, I608=>output_MAC_2_608, I609=>output_MAC_2_609, I610=>output_MAC_2_610, I611=>output_MAC_2_611, I612=>output_MAC_2_612, I613=>output_MAC_2_613, I614=>output_MAC_2_614, I615=>output_MAC_2_615, I616=>output_MAC_2_616, I617=>output_MAC_2_617, I618=>output_MAC_2_618, I619=>output_MAC_2_619, I620=>output_MAC_2_620, I621=>output_MAC_2_621, I622=>output_MAC_2_622, I623=>output_MAC_2_623, I624=>output_MAC_2_624, I625=>output_MAC_2_625, I626=>output_MAC_2_626, I627=>output_MAC_2_627, I628=>output_MAC_2_628, I629=>output_MAC_2_629, I630=>output_MAC_2_630, I631=>output_MAC_2_631, I632=>output_MAC_2_632, I633=>output_MAC_2_633, I634=>output_MAC_2_634, I635=>output_MAC_2_635, I636=>output_MAC_2_636, I637=>output_MAC_2_637, I638=>output_MAC_2_638, I639=>output_MAC_2_639, I640=>output_MAC_2_640, I641=>output_MAC_2_641, I642=>output_MAC_2_642, I643=>output_MAC_2_643, I644=>output_MAC_2_644, I645=>output_MAC_2_645, I646=>output_MAC_2_646, I647=>output_MAC_2_647, I648=>output_MAC_2_648, I649=>output_MAC_2_649, I650=>output_MAC_2_650, I651=>output_MAC_2_651, I652=>output_MAC_2_652, I653=>output_MAC_2_653, I654=>output_MAC_2_654, I655=>output_MAC_2_655, I656=>output_MAC_2_656, I657=>output_MAC_2_657, I658=>output_MAC_2_658, I659=>output_MAC_2_659, I660=>output_MAC_2_660, I661=>output_MAC_2_661, I662=>output_MAC_2_662, I663=>output_MAC_2_663, I664=>output_MAC_2_664, I665=>output_MAC_2_665, I666=>output_MAC_2_666, I667=>output_MAC_2_667, I668=>output_MAC_2_668, I669=>output_MAC_2_669, I670=>output_MAC_2_670, I671=>output_MAC_2_671, I672=>output_MAC_2_672, I673=>output_MAC_2_673, I674=>output_MAC_2_674, I675=>output_MAC_2_675, I676=>output_MAC_2_676, I677=>output_MAC_2_677, I678=>output_MAC_2_678, I679=>output_MAC_2_679, I680=>output_MAC_2_680, I681=>output_MAC_2_681, I682=>output_MAC_2_682, I683=>output_MAC_2_683, I684=>output_MAC_2_684, I685=>output_MAC_2_685, I686=>output_MAC_2_686, I687=>output_MAC_2_687, I688=>output_MAC_2_688, I689=>output_MAC_2_689, I690=>output_MAC_2_690, I691=>output_MAC_2_691, I692=>output_MAC_2_692, I693=>output_MAC_2_693, I694=>output_MAC_2_694, I695=>output_MAC_2_695, I696=>output_MAC_2_696, I697=>output_MAC_2_697, I698=>output_MAC_2_698, I699=>output_MAC_2_699, I700=>output_MAC_2_700, I701=>output_MAC_2_701, I702=>output_MAC_2_702, I703=>output_MAC_2_703, I704=>output_MAC_2_704, I705=>output_MAC_2_705, I706=>output_MAC_2_706, I707=>output_MAC_2_707, I708=>output_MAC_2_708, I709=>output_MAC_2_709, I710=>output_MAC_2_710, I711=>output_MAC_2_711, I712=>output_MAC_2_712, I713=>output_MAC_2_713, I714=>output_MAC_2_714, I715=>output_MAC_2_715, I716=>output_MAC_2_716, I717=>output_MAC_2_717, I718=>output_MAC_2_718, I719=>output_MAC_2_719, I720=>output_MAC_2_720, I721=>output_MAC_2_721, I722=>output_MAC_2_722, I723=>output_MAC_2_723, I724=>output_MAC_2_724, I725=>output_MAC_2_725, I726=>output_MAC_2_726, I727=>output_MAC_2_727, I728=>output_MAC_2_728, I729=>output_MAC_2_729, I730=>output_MAC_2_730, I731=>output_MAC_2_731, I732=>output_MAC_2_732, I733=>output_MAC_2_733, I734=>output_MAC_2_734, I735=>output_MAC_2_735, I736=>output_MAC_2_736, I737=>output_MAC_2_737, I738=>output_MAC_2_738, I739=>output_MAC_2_739, I740=>output_MAC_2_740, I741=>output_MAC_2_741, I742=>output_MAC_2_742, I743=>output_MAC_2_743, I744=>output_MAC_2_744, I745=>output_MAC_2_745, I746=>output_MAC_2_746, I747=>output_MAC_2_747, I748=>output_MAC_2_748, I749=>output_MAC_2_749, I750=>output_MAC_2_750, I751=>output_MAC_2_751, I752=>output_MAC_2_752, I753=>output_MAC_2_753, I754=>output_MAC_2_754, I755=>output_MAC_2_755, I756=>output_MAC_2_756, I757=>output_MAC_2_757, I758=>output_MAC_2_758, I759=>output_MAC_2_759, I760=>output_MAC_2_760, I761=>output_MAC_2_761, I762=>output_MAC_2_762, I763=>output_MAC_2_763, I764=>output_MAC_2_764, I765=>output_MAC_2_765, I766=>output_MAC_2_766, I767=>output_MAC_2_767, 
		SEL_mux=>SEL_mux, O=>output_row_2);

	mux_row_3: mux_768to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_3_0, I1=>output_MAC_3_1, I2=>output_MAC_3_2, I3=>output_MAC_3_3, I4=>output_MAC_3_4, I5=>output_MAC_3_5, I6=>output_MAC_3_6, I7=>output_MAC_3_7, I8=>output_MAC_3_8, I9=>output_MAC_3_9, I10=>output_MAC_3_10, I11=>output_MAC_3_11, I12=>output_MAC_3_12, I13=>output_MAC_3_13, I14=>output_MAC_3_14, I15=>output_MAC_3_15, I16=>output_MAC_3_16, I17=>output_MAC_3_17, I18=>output_MAC_3_18, I19=>output_MAC_3_19, I20=>output_MAC_3_20, I21=>output_MAC_3_21, I22=>output_MAC_3_22, I23=>output_MAC_3_23, I24=>output_MAC_3_24, I25=>output_MAC_3_25, I26=>output_MAC_3_26, I27=>output_MAC_3_27, I28=>output_MAC_3_28, I29=>output_MAC_3_29, I30=>output_MAC_3_30, I31=>output_MAC_3_31, I32=>output_MAC_3_32, I33=>output_MAC_3_33, I34=>output_MAC_3_34, I35=>output_MAC_3_35, I36=>output_MAC_3_36, I37=>output_MAC_3_37, I38=>output_MAC_3_38, I39=>output_MAC_3_39, I40=>output_MAC_3_40, I41=>output_MAC_3_41, I42=>output_MAC_3_42, I43=>output_MAC_3_43, I44=>output_MAC_3_44, I45=>output_MAC_3_45, I46=>output_MAC_3_46, I47=>output_MAC_3_47, I48=>output_MAC_3_48, I49=>output_MAC_3_49, I50=>output_MAC_3_50, I51=>output_MAC_3_51, I52=>output_MAC_3_52, I53=>output_MAC_3_53, I54=>output_MAC_3_54, I55=>output_MAC_3_55, I56=>output_MAC_3_56, I57=>output_MAC_3_57, I58=>output_MAC_3_58, I59=>output_MAC_3_59, I60=>output_MAC_3_60, I61=>output_MAC_3_61, I62=>output_MAC_3_62, I63=>output_MAC_3_63, I64=>output_MAC_3_64, I65=>output_MAC_3_65, I66=>output_MAC_3_66, I67=>output_MAC_3_67, I68=>output_MAC_3_68, I69=>output_MAC_3_69, I70=>output_MAC_3_70, I71=>output_MAC_3_71, I72=>output_MAC_3_72, I73=>output_MAC_3_73, I74=>output_MAC_3_74, I75=>output_MAC_3_75, I76=>output_MAC_3_76, I77=>output_MAC_3_77, I78=>output_MAC_3_78, I79=>output_MAC_3_79, I80=>output_MAC_3_80, I81=>output_MAC_3_81, I82=>output_MAC_3_82, I83=>output_MAC_3_83, I84=>output_MAC_3_84, I85=>output_MAC_3_85, I86=>output_MAC_3_86, I87=>output_MAC_3_87, I88=>output_MAC_3_88, I89=>output_MAC_3_89, I90=>output_MAC_3_90, I91=>output_MAC_3_91, I92=>output_MAC_3_92, I93=>output_MAC_3_93, I94=>output_MAC_3_94, I95=>output_MAC_3_95, I96=>output_MAC_3_96, I97=>output_MAC_3_97, I98=>output_MAC_3_98, I99=>output_MAC_3_99, I100=>output_MAC_3_100, I101=>output_MAC_3_101, I102=>output_MAC_3_102, I103=>output_MAC_3_103, I104=>output_MAC_3_104, I105=>output_MAC_3_105, I106=>output_MAC_3_106, I107=>output_MAC_3_107, I108=>output_MAC_3_108, I109=>output_MAC_3_109, I110=>output_MAC_3_110, I111=>output_MAC_3_111, I112=>output_MAC_3_112, I113=>output_MAC_3_113, I114=>output_MAC_3_114, I115=>output_MAC_3_115, I116=>output_MAC_3_116, I117=>output_MAC_3_117, I118=>output_MAC_3_118, I119=>output_MAC_3_119, I120=>output_MAC_3_120, I121=>output_MAC_3_121, I122=>output_MAC_3_122, I123=>output_MAC_3_123, I124=>output_MAC_3_124, I125=>output_MAC_3_125, I126=>output_MAC_3_126, I127=>output_MAC_3_127, I128=>output_MAC_3_128, I129=>output_MAC_3_129, I130=>output_MAC_3_130, I131=>output_MAC_3_131, I132=>output_MAC_3_132, I133=>output_MAC_3_133, I134=>output_MAC_3_134, I135=>output_MAC_3_135, I136=>output_MAC_3_136, I137=>output_MAC_3_137, I138=>output_MAC_3_138, I139=>output_MAC_3_139, I140=>output_MAC_3_140, I141=>output_MAC_3_141, I142=>output_MAC_3_142, I143=>output_MAC_3_143, I144=>output_MAC_3_144, I145=>output_MAC_3_145, I146=>output_MAC_3_146, I147=>output_MAC_3_147, I148=>output_MAC_3_148, I149=>output_MAC_3_149, I150=>output_MAC_3_150, I151=>output_MAC_3_151, I152=>output_MAC_3_152, I153=>output_MAC_3_153, I154=>output_MAC_3_154, I155=>output_MAC_3_155, I156=>output_MAC_3_156, I157=>output_MAC_3_157, I158=>output_MAC_3_158, I159=>output_MAC_3_159, I160=>output_MAC_3_160, I161=>output_MAC_3_161, I162=>output_MAC_3_162, I163=>output_MAC_3_163, I164=>output_MAC_3_164, I165=>output_MAC_3_165, I166=>output_MAC_3_166, I167=>output_MAC_3_167, I168=>output_MAC_3_168, I169=>output_MAC_3_169, I170=>output_MAC_3_170, I171=>output_MAC_3_171, I172=>output_MAC_3_172, I173=>output_MAC_3_173, I174=>output_MAC_3_174, I175=>output_MAC_3_175, I176=>output_MAC_3_176, I177=>output_MAC_3_177, I178=>output_MAC_3_178, I179=>output_MAC_3_179, I180=>output_MAC_3_180, I181=>output_MAC_3_181, I182=>output_MAC_3_182, I183=>output_MAC_3_183, I184=>output_MAC_3_184, I185=>output_MAC_3_185, I186=>output_MAC_3_186, I187=>output_MAC_3_187, I188=>output_MAC_3_188, I189=>output_MAC_3_189, I190=>output_MAC_3_190, I191=>output_MAC_3_191, I192=>output_MAC_3_192, I193=>output_MAC_3_193, I194=>output_MAC_3_194, I195=>output_MAC_3_195, I196=>output_MAC_3_196, I197=>output_MAC_3_197, I198=>output_MAC_3_198, I199=>output_MAC_3_199, I200=>output_MAC_3_200, I201=>output_MAC_3_201, I202=>output_MAC_3_202, I203=>output_MAC_3_203, I204=>output_MAC_3_204, I205=>output_MAC_3_205, I206=>output_MAC_3_206, I207=>output_MAC_3_207, I208=>output_MAC_3_208, I209=>output_MAC_3_209, I210=>output_MAC_3_210, I211=>output_MAC_3_211, I212=>output_MAC_3_212, I213=>output_MAC_3_213, I214=>output_MAC_3_214, I215=>output_MAC_3_215, I216=>output_MAC_3_216, I217=>output_MAC_3_217, I218=>output_MAC_3_218, I219=>output_MAC_3_219, I220=>output_MAC_3_220, I221=>output_MAC_3_221, I222=>output_MAC_3_222, I223=>output_MAC_3_223, I224=>output_MAC_3_224, I225=>output_MAC_3_225, I226=>output_MAC_3_226, I227=>output_MAC_3_227, I228=>output_MAC_3_228, I229=>output_MAC_3_229, I230=>output_MAC_3_230, I231=>output_MAC_3_231, I232=>output_MAC_3_232, I233=>output_MAC_3_233, I234=>output_MAC_3_234, I235=>output_MAC_3_235, I236=>output_MAC_3_236, I237=>output_MAC_3_237, I238=>output_MAC_3_238, I239=>output_MAC_3_239, I240=>output_MAC_3_240, I241=>output_MAC_3_241, I242=>output_MAC_3_242, I243=>output_MAC_3_243, I244=>output_MAC_3_244, I245=>output_MAC_3_245, I246=>output_MAC_3_246, I247=>output_MAC_3_247, I248=>output_MAC_3_248, I249=>output_MAC_3_249, I250=>output_MAC_3_250, I251=>output_MAC_3_251, I252=>output_MAC_3_252, I253=>output_MAC_3_253, I254=>output_MAC_3_254, I255=>output_MAC_3_255, I256=>output_MAC_3_256, I257=>output_MAC_3_257, I258=>output_MAC_3_258, I259=>output_MAC_3_259, I260=>output_MAC_3_260, I261=>output_MAC_3_261, I262=>output_MAC_3_262, I263=>output_MAC_3_263, I264=>output_MAC_3_264, I265=>output_MAC_3_265, I266=>output_MAC_3_266, I267=>output_MAC_3_267, I268=>output_MAC_3_268, I269=>output_MAC_3_269, I270=>output_MAC_3_270, I271=>output_MAC_3_271, I272=>output_MAC_3_272, I273=>output_MAC_3_273, I274=>output_MAC_3_274, I275=>output_MAC_3_275, I276=>output_MAC_3_276, I277=>output_MAC_3_277, I278=>output_MAC_3_278, I279=>output_MAC_3_279, I280=>output_MAC_3_280, I281=>output_MAC_3_281, I282=>output_MAC_3_282, I283=>output_MAC_3_283, I284=>output_MAC_3_284, I285=>output_MAC_3_285, I286=>output_MAC_3_286, I287=>output_MAC_3_287, I288=>output_MAC_3_288, I289=>output_MAC_3_289, I290=>output_MAC_3_290, I291=>output_MAC_3_291, I292=>output_MAC_3_292, I293=>output_MAC_3_293, I294=>output_MAC_3_294, I295=>output_MAC_3_295, I296=>output_MAC_3_296, I297=>output_MAC_3_297, I298=>output_MAC_3_298, I299=>output_MAC_3_299, I300=>output_MAC_3_300, I301=>output_MAC_3_301, I302=>output_MAC_3_302, I303=>output_MAC_3_303, I304=>output_MAC_3_304, I305=>output_MAC_3_305, I306=>output_MAC_3_306, I307=>output_MAC_3_307, I308=>output_MAC_3_308, I309=>output_MAC_3_309, I310=>output_MAC_3_310, I311=>output_MAC_3_311, I312=>output_MAC_3_312, I313=>output_MAC_3_313, I314=>output_MAC_3_314, I315=>output_MAC_3_315, I316=>output_MAC_3_316, I317=>output_MAC_3_317, I318=>output_MAC_3_318, I319=>output_MAC_3_319, I320=>output_MAC_3_320, I321=>output_MAC_3_321, I322=>output_MAC_3_322, I323=>output_MAC_3_323, I324=>output_MAC_3_324, I325=>output_MAC_3_325, I326=>output_MAC_3_326, I327=>output_MAC_3_327, I328=>output_MAC_3_328, I329=>output_MAC_3_329, I330=>output_MAC_3_330, I331=>output_MAC_3_331, I332=>output_MAC_3_332, I333=>output_MAC_3_333, I334=>output_MAC_3_334, I335=>output_MAC_3_335, I336=>output_MAC_3_336, I337=>output_MAC_3_337, I338=>output_MAC_3_338, I339=>output_MAC_3_339, I340=>output_MAC_3_340, I341=>output_MAC_3_341, I342=>output_MAC_3_342, I343=>output_MAC_3_343, I344=>output_MAC_3_344, I345=>output_MAC_3_345, I346=>output_MAC_3_346, I347=>output_MAC_3_347, I348=>output_MAC_3_348, I349=>output_MAC_3_349, I350=>output_MAC_3_350, I351=>output_MAC_3_351, I352=>output_MAC_3_352, I353=>output_MAC_3_353, I354=>output_MAC_3_354, I355=>output_MAC_3_355, I356=>output_MAC_3_356, I357=>output_MAC_3_357, I358=>output_MAC_3_358, I359=>output_MAC_3_359, I360=>output_MAC_3_360, I361=>output_MAC_3_361, I362=>output_MAC_3_362, I363=>output_MAC_3_363, I364=>output_MAC_3_364, I365=>output_MAC_3_365, I366=>output_MAC_3_366, I367=>output_MAC_3_367, I368=>output_MAC_3_368, I369=>output_MAC_3_369, I370=>output_MAC_3_370, I371=>output_MAC_3_371, I372=>output_MAC_3_372, I373=>output_MAC_3_373, I374=>output_MAC_3_374, I375=>output_MAC_3_375, I376=>output_MAC_3_376, I377=>output_MAC_3_377, I378=>output_MAC_3_378, I379=>output_MAC_3_379, I380=>output_MAC_3_380, I381=>output_MAC_3_381, I382=>output_MAC_3_382, I383=>output_MAC_3_383, I384=>output_MAC_3_384, I385=>output_MAC_3_385, I386=>output_MAC_3_386, I387=>output_MAC_3_387, I388=>output_MAC_3_388, I389=>output_MAC_3_389, I390=>output_MAC_3_390, I391=>output_MAC_3_391, I392=>output_MAC_3_392, I393=>output_MAC_3_393, I394=>output_MAC_3_394, I395=>output_MAC_3_395, I396=>output_MAC_3_396, I397=>output_MAC_3_397, I398=>output_MAC_3_398, I399=>output_MAC_3_399, I400=>output_MAC_3_400, I401=>output_MAC_3_401, I402=>output_MAC_3_402, I403=>output_MAC_3_403, I404=>output_MAC_3_404, I405=>output_MAC_3_405, I406=>output_MAC_3_406, I407=>output_MAC_3_407, I408=>output_MAC_3_408, I409=>output_MAC_3_409, I410=>output_MAC_3_410, I411=>output_MAC_3_411, I412=>output_MAC_3_412, I413=>output_MAC_3_413, I414=>output_MAC_3_414, I415=>output_MAC_3_415, I416=>output_MAC_3_416, I417=>output_MAC_3_417, I418=>output_MAC_3_418, I419=>output_MAC_3_419, I420=>output_MAC_3_420, I421=>output_MAC_3_421, I422=>output_MAC_3_422, I423=>output_MAC_3_423, I424=>output_MAC_3_424, I425=>output_MAC_3_425, I426=>output_MAC_3_426, I427=>output_MAC_3_427, I428=>output_MAC_3_428, I429=>output_MAC_3_429, I430=>output_MAC_3_430, I431=>output_MAC_3_431, I432=>output_MAC_3_432, I433=>output_MAC_3_433, I434=>output_MAC_3_434, I435=>output_MAC_3_435, I436=>output_MAC_3_436, I437=>output_MAC_3_437, I438=>output_MAC_3_438, I439=>output_MAC_3_439, I440=>output_MAC_3_440, I441=>output_MAC_3_441, I442=>output_MAC_3_442, I443=>output_MAC_3_443, I444=>output_MAC_3_444, I445=>output_MAC_3_445, I446=>output_MAC_3_446, I447=>output_MAC_3_447, I448=>output_MAC_3_448, I449=>output_MAC_3_449, I450=>output_MAC_3_450, I451=>output_MAC_3_451, I452=>output_MAC_3_452, I453=>output_MAC_3_453, I454=>output_MAC_3_454, I455=>output_MAC_3_455, I456=>output_MAC_3_456, I457=>output_MAC_3_457, I458=>output_MAC_3_458, I459=>output_MAC_3_459, I460=>output_MAC_3_460, I461=>output_MAC_3_461, I462=>output_MAC_3_462, I463=>output_MAC_3_463, I464=>output_MAC_3_464, I465=>output_MAC_3_465, I466=>output_MAC_3_466, I467=>output_MAC_3_467, I468=>output_MAC_3_468, I469=>output_MAC_3_469, I470=>output_MAC_3_470, I471=>output_MAC_3_471, I472=>output_MAC_3_472, I473=>output_MAC_3_473, I474=>output_MAC_3_474, I475=>output_MAC_3_475, I476=>output_MAC_3_476, I477=>output_MAC_3_477, I478=>output_MAC_3_478, I479=>output_MAC_3_479, I480=>output_MAC_3_480, I481=>output_MAC_3_481, I482=>output_MAC_3_482, I483=>output_MAC_3_483, I484=>output_MAC_3_484, I485=>output_MAC_3_485, I486=>output_MAC_3_486, I487=>output_MAC_3_487, I488=>output_MAC_3_488, I489=>output_MAC_3_489, I490=>output_MAC_3_490, I491=>output_MAC_3_491, I492=>output_MAC_3_492, I493=>output_MAC_3_493, I494=>output_MAC_3_494, I495=>output_MAC_3_495, I496=>output_MAC_3_496, I497=>output_MAC_3_497, I498=>output_MAC_3_498, I499=>output_MAC_3_499, I500=>output_MAC_3_500, I501=>output_MAC_3_501, I502=>output_MAC_3_502, I503=>output_MAC_3_503, I504=>output_MAC_3_504, I505=>output_MAC_3_505, I506=>output_MAC_3_506, I507=>output_MAC_3_507, I508=>output_MAC_3_508, I509=>output_MAC_3_509, I510=>output_MAC_3_510, I511=>output_MAC_3_511, I512=>output_MAC_3_512, I513=>output_MAC_3_513, I514=>output_MAC_3_514, I515=>output_MAC_3_515, I516=>output_MAC_3_516, I517=>output_MAC_3_517, I518=>output_MAC_3_518, I519=>output_MAC_3_519, I520=>output_MAC_3_520, I521=>output_MAC_3_521, I522=>output_MAC_3_522, I523=>output_MAC_3_523, I524=>output_MAC_3_524, I525=>output_MAC_3_525, I526=>output_MAC_3_526, I527=>output_MAC_3_527, I528=>output_MAC_3_528, I529=>output_MAC_3_529, I530=>output_MAC_3_530, I531=>output_MAC_3_531, I532=>output_MAC_3_532, I533=>output_MAC_3_533, I534=>output_MAC_3_534, I535=>output_MAC_3_535, I536=>output_MAC_3_536, I537=>output_MAC_3_537, I538=>output_MAC_3_538, I539=>output_MAC_3_539, I540=>output_MAC_3_540, I541=>output_MAC_3_541, I542=>output_MAC_3_542, I543=>output_MAC_3_543, I544=>output_MAC_3_544, I545=>output_MAC_3_545, I546=>output_MAC_3_546, I547=>output_MAC_3_547, I548=>output_MAC_3_548, I549=>output_MAC_3_549, I550=>output_MAC_3_550, I551=>output_MAC_3_551, I552=>output_MAC_3_552, I553=>output_MAC_3_553, I554=>output_MAC_3_554, I555=>output_MAC_3_555, I556=>output_MAC_3_556, I557=>output_MAC_3_557, I558=>output_MAC_3_558, I559=>output_MAC_3_559, I560=>output_MAC_3_560, I561=>output_MAC_3_561, I562=>output_MAC_3_562, I563=>output_MAC_3_563, I564=>output_MAC_3_564, I565=>output_MAC_3_565, I566=>output_MAC_3_566, I567=>output_MAC_3_567, I568=>output_MAC_3_568, I569=>output_MAC_3_569, I570=>output_MAC_3_570, I571=>output_MAC_3_571, I572=>output_MAC_3_572, I573=>output_MAC_3_573, I574=>output_MAC_3_574, I575=>output_MAC_3_575, I576=>output_MAC_3_576, I577=>output_MAC_3_577, I578=>output_MAC_3_578, I579=>output_MAC_3_579, I580=>output_MAC_3_580, I581=>output_MAC_3_581, I582=>output_MAC_3_582, I583=>output_MAC_3_583, I584=>output_MAC_3_584, I585=>output_MAC_3_585, I586=>output_MAC_3_586, I587=>output_MAC_3_587, I588=>output_MAC_3_588, I589=>output_MAC_3_589, I590=>output_MAC_3_590, I591=>output_MAC_3_591, I592=>output_MAC_3_592, I593=>output_MAC_3_593, I594=>output_MAC_3_594, I595=>output_MAC_3_595, I596=>output_MAC_3_596, I597=>output_MAC_3_597, I598=>output_MAC_3_598, I599=>output_MAC_3_599, I600=>output_MAC_3_600, I601=>output_MAC_3_601, I602=>output_MAC_3_602, I603=>output_MAC_3_603, I604=>output_MAC_3_604, I605=>output_MAC_3_605, I606=>output_MAC_3_606, I607=>output_MAC_3_607, I608=>output_MAC_3_608, I609=>output_MAC_3_609, I610=>output_MAC_3_610, I611=>output_MAC_3_611, I612=>output_MAC_3_612, I613=>output_MAC_3_613, I614=>output_MAC_3_614, I615=>output_MAC_3_615, I616=>output_MAC_3_616, I617=>output_MAC_3_617, I618=>output_MAC_3_618, I619=>output_MAC_3_619, I620=>output_MAC_3_620, I621=>output_MAC_3_621, I622=>output_MAC_3_622, I623=>output_MAC_3_623, I624=>output_MAC_3_624, I625=>output_MAC_3_625, I626=>output_MAC_3_626, I627=>output_MAC_3_627, I628=>output_MAC_3_628, I629=>output_MAC_3_629, I630=>output_MAC_3_630, I631=>output_MAC_3_631, I632=>output_MAC_3_632, I633=>output_MAC_3_633, I634=>output_MAC_3_634, I635=>output_MAC_3_635, I636=>output_MAC_3_636, I637=>output_MAC_3_637, I638=>output_MAC_3_638, I639=>output_MAC_3_639, I640=>output_MAC_3_640, I641=>output_MAC_3_641, I642=>output_MAC_3_642, I643=>output_MAC_3_643, I644=>output_MAC_3_644, I645=>output_MAC_3_645, I646=>output_MAC_3_646, I647=>output_MAC_3_647, I648=>output_MAC_3_648, I649=>output_MAC_3_649, I650=>output_MAC_3_650, I651=>output_MAC_3_651, I652=>output_MAC_3_652, I653=>output_MAC_3_653, I654=>output_MAC_3_654, I655=>output_MAC_3_655, I656=>output_MAC_3_656, I657=>output_MAC_3_657, I658=>output_MAC_3_658, I659=>output_MAC_3_659, I660=>output_MAC_3_660, I661=>output_MAC_3_661, I662=>output_MAC_3_662, I663=>output_MAC_3_663, I664=>output_MAC_3_664, I665=>output_MAC_3_665, I666=>output_MAC_3_666, I667=>output_MAC_3_667, I668=>output_MAC_3_668, I669=>output_MAC_3_669, I670=>output_MAC_3_670, I671=>output_MAC_3_671, I672=>output_MAC_3_672, I673=>output_MAC_3_673, I674=>output_MAC_3_674, I675=>output_MAC_3_675, I676=>output_MAC_3_676, I677=>output_MAC_3_677, I678=>output_MAC_3_678, I679=>output_MAC_3_679, I680=>output_MAC_3_680, I681=>output_MAC_3_681, I682=>output_MAC_3_682, I683=>output_MAC_3_683, I684=>output_MAC_3_684, I685=>output_MAC_3_685, I686=>output_MAC_3_686, I687=>output_MAC_3_687, I688=>output_MAC_3_688, I689=>output_MAC_3_689, I690=>output_MAC_3_690, I691=>output_MAC_3_691, I692=>output_MAC_3_692, I693=>output_MAC_3_693, I694=>output_MAC_3_694, I695=>output_MAC_3_695, I696=>output_MAC_3_696, I697=>output_MAC_3_697, I698=>output_MAC_3_698, I699=>output_MAC_3_699, I700=>output_MAC_3_700, I701=>output_MAC_3_701, I702=>output_MAC_3_702, I703=>output_MAC_3_703, I704=>output_MAC_3_704, I705=>output_MAC_3_705, I706=>output_MAC_3_706, I707=>output_MAC_3_707, I708=>output_MAC_3_708, I709=>output_MAC_3_709, I710=>output_MAC_3_710, I711=>output_MAC_3_711, I712=>output_MAC_3_712, I713=>output_MAC_3_713, I714=>output_MAC_3_714, I715=>output_MAC_3_715, I716=>output_MAC_3_716, I717=>output_MAC_3_717, I718=>output_MAC_3_718, I719=>output_MAC_3_719, I720=>output_MAC_3_720, I721=>output_MAC_3_721, I722=>output_MAC_3_722, I723=>output_MAC_3_723, I724=>output_MAC_3_724, I725=>output_MAC_3_725, I726=>output_MAC_3_726, I727=>output_MAC_3_727, I728=>output_MAC_3_728, I729=>output_MAC_3_729, I730=>output_MAC_3_730, I731=>output_MAC_3_731, I732=>output_MAC_3_732, I733=>output_MAC_3_733, I734=>output_MAC_3_734, I735=>output_MAC_3_735, I736=>output_MAC_3_736, I737=>output_MAC_3_737, I738=>output_MAC_3_738, I739=>output_MAC_3_739, I740=>output_MAC_3_740, I741=>output_MAC_3_741, I742=>output_MAC_3_742, I743=>output_MAC_3_743, I744=>output_MAC_3_744, I745=>output_MAC_3_745, I746=>output_MAC_3_746, I747=>output_MAC_3_747, I748=>output_MAC_3_748, I749=>output_MAC_3_749, I750=>output_MAC_3_750, I751=>output_MAC_3_751, I752=>output_MAC_3_752, I753=>output_MAC_3_753, I754=>output_MAC_3_754, I755=>output_MAC_3_755, I756=>output_MAC_3_756, I757=>output_MAC_3_757, I758=>output_MAC_3_758, I759=>output_MAC_3_759, I760=>output_MAC_3_760, I761=>output_MAC_3_761, I762=>output_MAC_3_762, I763=>output_MAC_3_763, I764=>output_MAC_3_764, I765=>output_MAC_3_765, I766=>output_MAC_3_766, I767=>output_MAC_3_767, 
		SEL_mux=>SEL_mux, O=>output_row_3);

	mux_row_4: mux_768to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_4_0, I1=>output_MAC_4_1, I2=>output_MAC_4_2, I3=>output_MAC_4_3, I4=>output_MAC_4_4, I5=>output_MAC_4_5, I6=>output_MAC_4_6, I7=>output_MAC_4_7, I8=>output_MAC_4_8, I9=>output_MAC_4_9, I10=>output_MAC_4_10, I11=>output_MAC_4_11, I12=>output_MAC_4_12, I13=>output_MAC_4_13, I14=>output_MAC_4_14, I15=>output_MAC_4_15, I16=>output_MAC_4_16, I17=>output_MAC_4_17, I18=>output_MAC_4_18, I19=>output_MAC_4_19, I20=>output_MAC_4_20, I21=>output_MAC_4_21, I22=>output_MAC_4_22, I23=>output_MAC_4_23, I24=>output_MAC_4_24, I25=>output_MAC_4_25, I26=>output_MAC_4_26, I27=>output_MAC_4_27, I28=>output_MAC_4_28, I29=>output_MAC_4_29, I30=>output_MAC_4_30, I31=>output_MAC_4_31, I32=>output_MAC_4_32, I33=>output_MAC_4_33, I34=>output_MAC_4_34, I35=>output_MAC_4_35, I36=>output_MAC_4_36, I37=>output_MAC_4_37, I38=>output_MAC_4_38, I39=>output_MAC_4_39, I40=>output_MAC_4_40, I41=>output_MAC_4_41, I42=>output_MAC_4_42, I43=>output_MAC_4_43, I44=>output_MAC_4_44, I45=>output_MAC_4_45, I46=>output_MAC_4_46, I47=>output_MAC_4_47, I48=>output_MAC_4_48, I49=>output_MAC_4_49, I50=>output_MAC_4_50, I51=>output_MAC_4_51, I52=>output_MAC_4_52, I53=>output_MAC_4_53, I54=>output_MAC_4_54, I55=>output_MAC_4_55, I56=>output_MAC_4_56, I57=>output_MAC_4_57, I58=>output_MAC_4_58, I59=>output_MAC_4_59, I60=>output_MAC_4_60, I61=>output_MAC_4_61, I62=>output_MAC_4_62, I63=>output_MAC_4_63, I64=>output_MAC_4_64, I65=>output_MAC_4_65, I66=>output_MAC_4_66, I67=>output_MAC_4_67, I68=>output_MAC_4_68, I69=>output_MAC_4_69, I70=>output_MAC_4_70, I71=>output_MAC_4_71, I72=>output_MAC_4_72, I73=>output_MAC_4_73, I74=>output_MAC_4_74, I75=>output_MAC_4_75, I76=>output_MAC_4_76, I77=>output_MAC_4_77, I78=>output_MAC_4_78, I79=>output_MAC_4_79, I80=>output_MAC_4_80, I81=>output_MAC_4_81, I82=>output_MAC_4_82, I83=>output_MAC_4_83, I84=>output_MAC_4_84, I85=>output_MAC_4_85, I86=>output_MAC_4_86, I87=>output_MAC_4_87, I88=>output_MAC_4_88, I89=>output_MAC_4_89, I90=>output_MAC_4_90, I91=>output_MAC_4_91, I92=>output_MAC_4_92, I93=>output_MAC_4_93, I94=>output_MAC_4_94, I95=>output_MAC_4_95, I96=>output_MAC_4_96, I97=>output_MAC_4_97, I98=>output_MAC_4_98, I99=>output_MAC_4_99, I100=>output_MAC_4_100, I101=>output_MAC_4_101, I102=>output_MAC_4_102, I103=>output_MAC_4_103, I104=>output_MAC_4_104, I105=>output_MAC_4_105, I106=>output_MAC_4_106, I107=>output_MAC_4_107, I108=>output_MAC_4_108, I109=>output_MAC_4_109, I110=>output_MAC_4_110, I111=>output_MAC_4_111, I112=>output_MAC_4_112, I113=>output_MAC_4_113, I114=>output_MAC_4_114, I115=>output_MAC_4_115, I116=>output_MAC_4_116, I117=>output_MAC_4_117, I118=>output_MAC_4_118, I119=>output_MAC_4_119, I120=>output_MAC_4_120, I121=>output_MAC_4_121, I122=>output_MAC_4_122, I123=>output_MAC_4_123, I124=>output_MAC_4_124, I125=>output_MAC_4_125, I126=>output_MAC_4_126, I127=>output_MAC_4_127, I128=>output_MAC_4_128, I129=>output_MAC_4_129, I130=>output_MAC_4_130, I131=>output_MAC_4_131, I132=>output_MAC_4_132, I133=>output_MAC_4_133, I134=>output_MAC_4_134, I135=>output_MAC_4_135, I136=>output_MAC_4_136, I137=>output_MAC_4_137, I138=>output_MAC_4_138, I139=>output_MAC_4_139, I140=>output_MAC_4_140, I141=>output_MAC_4_141, I142=>output_MAC_4_142, I143=>output_MAC_4_143, I144=>output_MAC_4_144, I145=>output_MAC_4_145, I146=>output_MAC_4_146, I147=>output_MAC_4_147, I148=>output_MAC_4_148, I149=>output_MAC_4_149, I150=>output_MAC_4_150, I151=>output_MAC_4_151, I152=>output_MAC_4_152, I153=>output_MAC_4_153, I154=>output_MAC_4_154, I155=>output_MAC_4_155, I156=>output_MAC_4_156, I157=>output_MAC_4_157, I158=>output_MAC_4_158, I159=>output_MAC_4_159, I160=>output_MAC_4_160, I161=>output_MAC_4_161, I162=>output_MAC_4_162, I163=>output_MAC_4_163, I164=>output_MAC_4_164, I165=>output_MAC_4_165, I166=>output_MAC_4_166, I167=>output_MAC_4_167, I168=>output_MAC_4_168, I169=>output_MAC_4_169, I170=>output_MAC_4_170, I171=>output_MAC_4_171, I172=>output_MAC_4_172, I173=>output_MAC_4_173, I174=>output_MAC_4_174, I175=>output_MAC_4_175, I176=>output_MAC_4_176, I177=>output_MAC_4_177, I178=>output_MAC_4_178, I179=>output_MAC_4_179, I180=>output_MAC_4_180, I181=>output_MAC_4_181, I182=>output_MAC_4_182, I183=>output_MAC_4_183, I184=>output_MAC_4_184, I185=>output_MAC_4_185, I186=>output_MAC_4_186, I187=>output_MAC_4_187, I188=>output_MAC_4_188, I189=>output_MAC_4_189, I190=>output_MAC_4_190, I191=>output_MAC_4_191, I192=>output_MAC_4_192, I193=>output_MAC_4_193, I194=>output_MAC_4_194, I195=>output_MAC_4_195, I196=>output_MAC_4_196, I197=>output_MAC_4_197, I198=>output_MAC_4_198, I199=>output_MAC_4_199, I200=>output_MAC_4_200, I201=>output_MAC_4_201, I202=>output_MAC_4_202, I203=>output_MAC_4_203, I204=>output_MAC_4_204, I205=>output_MAC_4_205, I206=>output_MAC_4_206, I207=>output_MAC_4_207, I208=>output_MAC_4_208, I209=>output_MAC_4_209, I210=>output_MAC_4_210, I211=>output_MAC_4_211, I212=>output_MAC_4_212, I213=>output_MAC_4_213, I214=>output_MAC_4_214, I215=>output_MAC_4_215, I216=>output_MAC_4_216, I217=>output_MAC_4_217, I218=>output_MAC_4_218, I219=>output_MAC_4_219, I220=>output_MAC_4_220, I221=>output_MAC_4_221, I222=>output_MAC_4_222, I223=>output_MAC_4_223, I224=>output_MAC_4_224, I225=>output_MAC_4_225, I226=>output_MAC_4_226, I227=>output_MAC_4_227, I228=>output_MAC_4_228, I229=>output_MAC_4_229, I230=>output_MAC_4_230, I231=>output_MAC_4_231, I232=>output_MAC_4_232, I233=>output_MAC_4_233, I234=>output_MAC_4_234, I235=>output_MAC_4_235, I236=>output_MAC_4_236, I237=>output_MAC_4_237, I238=>output_MAC_4_238, I239=>output_MAC_4_239, I240=>output_MAC_4_240, I241=>output_MAC_4_241, I242=>output_MAC_4_242, I243=>output_MAC_4_243, I244=>output_MAC_4_244, I245=>output_MAC_4_245, I246=>output_MAC_4_246, I247=>output_MAC_4_247, I248=>output_MAC_4_248, I249=>output_MAC_4_249, I250=>output_MAC_4_250, I251=>output_MAC_4_251, I252=>output_MAC_4_252, I253=>output_MAC_4_253, I254=>output_MAC_4_254, I255=>output_MAC_4_255, I256=>output_MAC_4_256, I257=>output_MAC_4_257, I258=>output_MAC_4_258, I259=>output_MAC_4_259, I260=>output_MAC_4_260, I261=>output_MAC_4_261, I262=>output_MAC_4_262, I263=>output_MAC_4_263, I264=>output_MAC_4_264, I265=>output_MAC_4_265, I266=>output_MAC_4_266, I267=>output_MAC_4_267, I268=>output_MAC_4_268, I269=>output_MAC_4_269, I270=>output_MAC_4_270, I271=>output_MAC_4_271, I272=>output_MAC_4_272, I273=>output_MAC_4_273, I274=>output_MAC_4_274, I275=>output_MAC_4_275, I276=>output_MAC_4_276, I277=>output_MAC_4_277, I278=>output_MAC_4_278, I279=>output_MAC_4_279, I280=>output_MAC_4_280, I281=>output_MAC_4_281, I282=>output_MAC_4_282, I283=>output_MAC_4_283, I284=>output_MAC_4_284, I285=>output_MAC_4_285, I286=>output_MAC_4_286, I287=>output_MAC_4_287, I288=>output_MAC_4_288, I289=>output_MAC_4_289, I290=>output_MAC_4_290, I291=>output_MAC_4_291, I292=>output_MAC_4_292, I293=>output_MAC_4_293, I294=>output_MAC_4_294, I295=>output_MAC_4_295, I296=>output_MAC_4_296, I297=>output_MAC_4_297, I298=>output_MAC_4_298, I299=>output_MAC_4_299, I300=>output_MAC_4_300, I301=>output_MAC_4_301, I302=>output_MAC_4_302, I303=>output_MAC_4_303, I304=>output_MAC_4_304, I305=>output_MAC_4_305, I306=>output_MAC_4_306, I307=>output_MAC_4_307, I308=>output_MAC_4_308, I309=>output_MAC_4_309, I310=>output_MAC_4_310, I311=>output_MAC_4_311, I312=>output_MAC_4_312, I313=>output_MAC_4_313, I314=>output_MAC_4_314, I315=>output_MAC_4_315, I316=>output_MAC_4_316, I317=>output_MAC_4_317, I318=>output_MAC_4_318, I319=>output_MAC_4_319, I320=>output_MAC_4_320, I321=>output_MAC_4_321, I322=>output_MAC_4_322, I323=>output_MAC_4_323, I324=>output_MAC_4_324, I325=>output_MAC_4_325, I326=>output_MAC_4_326, I327=>output_MAC_4_327, I328=>output_MAC_4_328, I329=>output_MAC_4_329, I330=>output_MAC_4_330, I331=>output_MAC_4_331, I332=>output_MAC_4_332, I333=>output_MAC_4_333, I334=>output_MAC_4_334, I335=>output_MAC_4_335, I336=>output_MAC_4_336, I337=>output_MAC_4_337, I338=>output_MAC_4_338, I339=>output_MAC_4_339, I340=>output_MAC_4_340, I341=>output_MAC_4_341, I342=>output_MAC_4_342, I343=>output_MAC_4_343, I344=>output_MAC_4_344, I345=>output_MAC_4_345, I346=>output_MAC_4_346, I347=>output_MAC_4_347, I348=>output_MAC_4_348, I349=>output_MAC_4_349, I350=>output_MAC_4_350, I351=>output_MAC_4_351, I352=>output_MAC_4_352, I353=>output_MAC_4_353, I354=>output_MAC_4_354, I355=>output_MAC_4_355, I356=>output_MAC_4_356, I357=>output_MAC_4_357, I358=>output_MAC_4_358, I359=>output_MAC_4_359, I360=>output_MAC_4_360, I361=>output_MAC_4_361, I362=>output_MAC_4_362, I363=>output_MAC_4_363, I364=>output_MAC_4_364, I365=>output_MAC_4_365, I366=>output_MAC_4_366, I367=>output_MAC_4_367, I368=>output_MAC_4_368, I369=>output_MAC_4_369, I370=>output_MAC_4_370, I371=>output_MAC_4_371, I372=>output_MAC_4_372, I373=>output_MAC_4_373, I374=>output_MAC_4_374, I375=>output_MAC_4_375, I376=>output_MAC_4_376, I377=>output_MAC_4_377, I378=>output_MAC_4_378, I379=>output_MAC_4_379, I380=>output_MAC_4_380, I381=>output_MAC_4_381, I382=>output_MAC_4_382, I383=>output_MAC_4_383, I384=>output_MAC_4_384, I385=>output_MAC_4_385, I386=>output_MAC_4_386, I387=>output_MAC_4_387, I388=>output_MAC_4_388, I389=>output_MAC_4_389, I390=>output_MAC_4_390, I391=>output_MAC_4_391, I392=>output_MAC_4_392, I393=>output_MAC_4_393, I394=>output_MAC_4_394, I395=>output_MAC_4_395, I396=>output_MAC_4_396, I397=>output_MAC_4_397, I398=>output_MAC_4_398, I399=>output_MAC_4_399, I400=>output_MAC_4_400, I401=>output_MAC_4_401, I402=>output_MAC_4_402, I403=>output_MAC_4_403, I404=>output_MAC_4_404, I405=>output_MAC_4_405, I406=>output_MAC_4_406, I407=>output_MAC_4_407, I408=>output_MAC_4_408, I409=>output_MAC_4_409, I410=>output_MAC_4_410, I411=>output_MAC_4_411, I412=>output_MAC_4_412, I413=>output_MAC_4_413, I414=>output_MAC_4_414, I415=>output_MAC_4_415, I416=>output_MAC_4_416, I417=>output_MAC_4_417, I418=>output_MAC_4_418, I419=>output_MAC_4_419, I420=>output_MAC_4_420, I421=>output_MAC_4_421, I422=>output_MAC_4_422, I423=>output_MAC_4_423, I424=>output_MAC_4_424, I425=>output_MAC_4_425, I426=>output_MAC_4_426, I427=>output_MAC_4_427, I428=>output_MAC_4_428, I429=>output_MAC_4_429, I430=>output_MAC_4_430, I431=>output_MAC_4_431, I432=>output_MAC_4_432, I433=>output_MAC_4_433, I434=>output_MAC_4_434, I435=>output_MAC_4_435, I436=>output_MAC_4_436, I437=>output_MAC_4_437, I438=>output_MAC_4_438, I439=>output_MAC_4_439, I440=>output_MAC_4_440, I441=>output_MAC_4_441, I442=>output_MAC_4_442, I443=>output_MAC_4_443, I444=>output_MAC_4_444, I445=>output_MAC_4_445, I446=>output_MAC_4_446, I447=>output_MAC_4_447, I448=>output_MAC_4_448, I449=>output_MAC_4_449, I450=>output_MAC_4_450, I451=>output_MAC_4_451, I452=>output_MAC_4_452, I453=>output_MAC_4_453, I454=>output_MAC_4_454, I455=>output_MAC_4_455, I456=>output_MAC_4_456, I457=>output_MAC_4_457, I458=>output_MAC_4_458, I459=>output_MAC_4_459, I460=>output_MAC_4_460, I461=>output_MAC_4_461, I462=>output_MAC_4_462, I463=>output_MAC_4_463, I464=>output_MAC_4_464, I465=>output_MAC_4_465, I466=>output_MAC_4_466, I467=>output_MAC_4_467, I468=>output_MAC_4_468, I469=>output_MAC_4_469, I470=>output_MAC_4_470, I471=>output_MAC_4_471, I472=>output_MAC_4_472, I473=>output_MAC_4_473, I474=>output_MAC_4_474, I475=>output_MAC_4_475, I476=>output_MAC_4_476, I477=>output_MAC_4_477, I478=>output_MAC_4_478, I479=>output_MAC_4_479, I480=>output_MAC_4_480, I481=>output_MAC_4_481, I482=>output_MAC_4_482, I483=>output_MAC_4_483, I484=>output_MAC_4_484, I485=>output_MAC_4_485, I486=>output_MAC_4_486, I487=>output_MAC_4_487, I488=>output_MAC_4_488, I489=>output_MAC_4_489, I490=>output_MAC_4_490, I491=>output_MAC_4_491, I492=>output_MAC_4_492, I493=>output_MAC_4_493, I494=>output_MAC_4_494, I495=>output_MAC_4_495, I496=>output_MAC_4_496, I497=>output_MAC_4_497, I498=>output_MAC_4_498, I499=>output_MAC_4_499, I500=>output_MAC_4_500, I501=>output_MAC_4_501, I502=>output_MAC_4_502, I503=>output_MAC_4_503, I504=>output_MAC_4_504, I505=>output_MAC_4_505, I506=>output_MAC_4_506, I507=>output_MAC_4_507, I508=>output_MAC_4_508, I509=>output_MAC_4_509, I510=>output_MAC_4_510, I511=>output_MAC_4_511, I512=>output_MAC_4_512, I513=>output_MAC_4_513, I514=>output_MAC_4_514, I515=>output_MAC_4_515, I516=>output_MAC_4_516, I517=>output_MAC_4_517, I518=>output_MAC_4_518, I519=>output_MAC_4_519, I520=>output_MAC_4_520, I521=>output_MAC_4_521, I522=>output_MAC_4_522, I523=>output_MAC_4_523, I524=>output_MAC_4_524, I525=>output_MAC_4_525, I526=>output_MAC_4_526, I527=>output_MAC_4_527, I528=>output_MAC_4_528, I529=>output_MAC_4_529, I530=>output_MAC_4_530, I531=>output_MAC_4_531, I532=>output_MAC_4_532, I533=>output_MAC_4_533, I534=>output_MAC_4_534, I535=>output_MAC_4_535, I536=>output_MAC_4_536, I537=>output_MAC_4_537, I538=>output_MAC_4_538, I539=>output_MAC_4_539, I540=>output_MAC_4_540, I541=>output_MAC_4_541, I542=>output_MAC_4_542, I543=>output_MAC_4_543, I544=>output_MAC_4_544, I545=>output_MAC_4_545, I546=>output_MAC_4_546, I547=>output_MAC_4_547, I548=>output_MAC_4_548, I549=>output_MAC_4_549, I550=>output_MAC_4_550, I551=>output_MAC_4_551, I552=>output_MAC_4_552, I553=>output_MAC_4_553, I554=>output_MAC_4_554, I555=>output_MAC_4_555, I556=>output_MAC_4_556, I557=>output_MAC_4_557, I558=>output_MAC_4_558, I559=>output_MAC_4_559, I560=>output_MAC_4_560, I561=>output_MAC_4_561, I562=>output_MAC_4_562, I563=>output_MAC_4_563, I564=>output_MAC_4_564, I565=>output_MAC_4_565, I566=>output_MAC_4_566, I567=>output_MAC_4_567, I568=>output_MAC_4_568, I569=>output_MAC_4_569, I570=>output_MAC_4_570, I571=>output_MAC_4_571, I572=>output_MAC_4_572, I573=>output_MAC_4_573, I574=>output_MAC_4_574, I575=>output_MAC_4_575, I576=>output_MAC_4_576, I577=>output_MAC_4_577, I578=>output_MAC_4_578, I579=>output_MAC_4_579, I580=>output_MAC_4_580, I581=>output_MAC_4_581, I582=>output_MAC_4_582, I583=>output_MAC_4_583, I584=>output_MAC_4_584, I585=>output_MAC_4_585, I586=>output_MAC_4_586, I587=>output_MAC_4_587, I588=>output_MAC_4_588, I589=>output_MAC_4_589, I590=>output_MAC_4_590, I591=>output_MAC_4_591, I592=>output_MAC_4_592, I593=>output_MAC_4_593, I594=>output_MAC_4_594, I595=>output_MAC_4_595, I596=>output_MAC_4_596, I597=>output_MAC_4_597, I598=>output_MAC_4_598, I599=>output_MAC_4_599, I600=>output_MAC_4_600, I601=>output_MAC_4_601, I602=>output_MAC_4_602, I603=>output_MAC_4_603, I604=>output_MAC_4_604, I605=>output_MAC_4_605, I606=>output_MAC_4_606, I607=>output_MAC_4_607, I608=>output_MAC_4_608, I609=>output_MAC_4_609, I610=>output_MAC_4_610, I611=>output_MAC_4_611, I612=>output_MAC_4_612, I613=>output_MAC_4_613, I614=>output_MAC_4_614, I615=>output_MAC_4_615, I616=>output_MAC_4_616, I617=>output_MAC_4_617, I618=>output_MAC_4_618, I619=>output_MAC_4_619, I620=>output_MAC_4_620, I621=>output_MAC_4_621, I622=>output_MAC_4_622, I623=>output_MAC_4_623, I624=>output_MAC_4_624, I625=>output_MAC_4_625, I626=>output_MAC_4_626, I627=>output_MAC_4_627, I628=>output_MAC_4_628, I629=>output_MAC_4_629, I630=>output_MAC_4_630, I631=>output_MAC_4_631, I632=>output_MAC_4_632, I633=>output_MAC_4_633, I634=>output_MAC_4_634, I635=>output_MAC_4_635, I636=>output_MAC_4_636, I637=>output_MAC_4_637, I638=>output_MAC_4_638, I639=>output_MAC_4_639, I640=>output_MAC_4_640, I641=>output_MAC_4_641, I642=>output_MAC_4_642, I643=>output_MAC_4_643, I644=>output_MAC_4_644, I645=>output_MAC_4_645, I646=>output_MAC_4_646, I647=>output_MAC_4_647, I648=>output_MAC_4_648, I649=>output_MAC_4_649, I650=>output_MAC_4_650, I651=>output_MAC_4_651, I652=>output_MAC_4_652, I653=>output_MAC_4_653, I654=>output_MAC_4_654, I655=>output_MAC_4_655, I656=>output_MAC_4_656, I657=>output_MAC_4_657, I658=>output_MAC_4_658, I659=>output_MAC_4_659, I660=>output_MAC_4_660, I661=>output_MAC_4_661, I662=>output_MAC_4_662, I663=>output_MAC_4_663, I664=>output_MAC_4_664, I665=>output_MAC_4_665, I666=>output_MAC_4_666, I667=>output_MAC_4_667, I668=>output_MAC_4_668, I669=>output_MAC_4_669, I670=>output_MAC_4_670, I671=>output_MAC_4_671, I672=>output_MAC_4_672, I673=>output_MAC_4_673, I674=>output_MAC_4_674, I675=>output_MAC_4_675, I676=>output_MAC_4_676, I677=>output_MAC_4_677, I678=>output_MAC_4_678, I679=>output_MAC_4_679, I680=>output_MAC_4_680, I681=>output_MAC_4_681, I682=>output_MAC_4_682, I683=>output_MAC_4_683, I684=>output_MAC_4_684, I685=>output_MAC_4_685, I686=>output_MAC_4_686, I687=>output_MAC_4_687, I688=>output_MAC_4_688, I689=>output_MAC_4_689, I690=>output_MAC_4_690, I691=>output_MAC_4_691, I692=>output_MAC_4_692, I693=>output_MAC_4_693, I694=>output_MAC_4_694, I695=>output_MAC_4_695, I696=>output_MAC_4_696, I697=>output_MAC_4_697, I698=>output_MAC_4_698, I699=>output_MAC_4_699, I700=>output_MAC_4_700, I701=>output_MAC_4_701, I702=>output_MAC_4_702, I703=>output_MAC_4_703, I704=>output_MAC_4_704, I705=>output_MAC_4_705, I706=>output_MAC_4_706, I707=>output_MAC_4_707, I708=>output_MAC_4_708, I709=>output_MAC_4_709, I710=>output_MAC_4_710, I711=>output_MAC_4_711, I712=>output_MAC_4_712, I713=>output_MAC_4_713, I714=>output_MAC_4_714, I715=>output_MAC_4_715, I716=>output_MAC_4_716, I717=>output_MAC_4_717, I718=>output_MAC_4_718, I719=>output_MAC_4_719, I720=>output_MAC_4_720, I721=>output_MAC_4_721, I722=>output_MAC_4_722, I723=>output_MAC_4_723, I724=>output_MAC_4_724, I725=>output_MAC_4_725, I726=>output_MAC_4_726, I727=>output_MAC_4_727, I728=>output_MAC_4_728, I729=>output_MAC_4_729, I730=>output_MAC_4_730, I731=>output_MAC_4_731, I732=>output_MAC_4_732, I733=>output_MAC_4_733, I734=>output_MAC_4_734, I735=>output_MAC_4_735, I736=>output_MAC_4_736, I737=>output_MAC_4_737, I738=>output_MAC_4_738, I739=>output_MAC_4_739, I740=>output_MAC_4_740, I741=>output_MAC_4_741, I742=>output_MAC_4_742, I743=>output_MAC_4_743, I744=>output_MAC_4_744, I745=>output_MAC_4_745, I746=>output_MAC_4_746, I747=>output_MAC_4_747, I748=>output_MAC_4_748, I749=>output_MAC_4_749, I750=>output_MAC_4_750, I751=>output_MAC_4_751, I752=>output_MAC_4_752, I753=>output_MAC_4_753, I754=>output_MAC_4_754, I755=>output_MAC_4_755, I756=>output_MAC_4_756, I757=>output_MAC_4_757, I758=>output_MAC_4_758, I759=>output_MAC_4_759, I760=>output_MAC_4_760, I761=>output_MAC_4_761, I762=>output_MAC_4_762, I763=>output_MAC_4_763, I764=>output_MAC_4_764, I765=>output_MAC_4_765, I766=>output_MAC_4_766, I767=>output_MAC_4_767, 
		SEL_mux=>SEL_mux, O=>output_row_4);

	mux_row_5: mux_768to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_5_0, I1=>output_MAC_5_1, I2=>output_MAC_5_2, I3=>output_MAC_5_3, I4=>output_MAC_5_4, I5=>output_MAC_5_5, I6=>output_MAC_5_6, I7=>output_MAC_5_7, I8=>output_MAC_5_8, I9=>output_MAC_5_9, I10=>output_MAC_5_10, I11=>output_MAC_5_11, I12=>output_MAC_5_12, I13=>output_MAC_5_13, I14=>output_MAC_5_14, I15=>output_MAC_5_15, I16=>output_MAC_5_16, I17=>output_MAC_5_17, I18=>output_MAC_5_18, I19=>output_MAC_5_19, I20=>output_MAC_5_20, I21=>output_MAC_5_21, I22=>output_MAC_5_22, I23=>output_MAC_5_23, I24=>output_MAC_5_24, I25=>output_MAC_5_25, I26=>output_MAC_5_26, I27=>output_MAC_5_27, I28=>output_MAC_5_28, I29=>output_MAC_5_29, I30=>output_MAC_5_30, I31=>output_MAC_5_31, I32=>output_MAC_5_32, I33=>output_MAC_5_33, I34=>output_MAC_5_34, I35=>output_MAC_5_35, I36=>output_MAC_5_36, I37=>output_MAC_5_37, I38=>output_MAC_5_38, I39=>output_MAC_5_39, I40=>output_MAC_5_40, I41=>output_MAC_5_41, I42=>output_MAC_5_42, I43=>output_MAC_5_43, I44=>output_MAC_5_44, I45=>output_MAC_5_45, I46=>output_MAC_5_46, I47=>output_MAC_5_47, I48=>output_MAC_5_48, I49=>output_MAC_5_49, I50=>output_MAC_5_50, I51=>output_MAC_5_51, I52=>output_MAC_5_52, I53=>output_MAC_5_53, I54=>output_MAC_5_54, I55=>output_MAC_5_55, I56=>output_MAC_5_56, I57=>output_MAC_5_57, I58=>output_MAC_5_58, I59=>output_MAC_5_59, I60=>output_MAC_5_60, I61=>output_MAC_5_61, I62=>output_MAC_5_62, I63=>output_MAC_5_63, I64=>output_MAC_5_64, I65=>output_MAC_5_65, I66=>output_MAC_5_66, I67=>output_MAC_5_67, I68=>output_MAC_5_68, I69=>output_MAC_5_69, I70=>output_MAC_5_70, I71=>output_MAC_5_71, I72=>output_MAC_5_72, I73=>output_MAC_5_73, I74=>output_MAC_5_74, I75=>output_MAC_5_75, I76=>output_MAC_5_76, I77=>output_MAC_5_77, I78=>output_MAC_5_78, I79=>output_MAC_5_79, I80=>output_MAC_5_80, I81=>output_MAC_5_81, I82=>output_MAC_5_82, I83=>output_MAC_5_83, I84=>output_MAC_5_84, I85=>output_MAC_5_85, I86=>output_MAC_5_86, I87=>output_MAC_5_87, I88=>output_MAC_5_88, I89=>output_MAC_5_89, I90=>output_MAC_5_90, I91=>output_MAC_5_91, I92=>output_MAC_5_92, I93=>output_MAC_5_93, I94=>output_MAC_5_94, I95=>output_MAC_5_95, I96=>output_MAC_5_96, I97=>output_MAC_5_97, I98=>output_MAC_5_98, I99=>output_MAC_5_99, I100=>output_MAC_5_100, I101=>output_MAC_5_101, I102=>output_MAC_5_102, I103=>output_MAC_5_103, I104=>output_MAC_5_104, I105=>output_MAC_5_105, I106=>output_MAC_5_106, I107=>output_MAC_5_107, I108=>output_MAC_5_108, I109=>output_MAC_5_109, I110=>output_MAC_5_110, I111=>output_MAC_5_111, I112=>output_MAC_5_112, I113=>output_MAC_5_113, I114=>output_MAC_5_114, I115=>output_MAC_5_115, I116=>output_MAC_5_116, I117=>output_MAC_5_117, I118=>output_MAC_5_118, I119=>output_MAC_5_119, I120=>output_MAC_5_120, I121=>output_MAC_5_121, I122=>output_MAC_5_122, I123=>output_MAC_5_123, I124=>output_MAC_5_124, I125=>output_MAC_5_125, I126=>output_MAC_5_126, I127=>output_MAC_5_127, I128=>output_MAC_5_128, I129=>output_MAC_5_129, I130=>output_MAC_5_130, I131=>output_MAC_5_131, I132=>output_MAC_5_132, I133=>output_MAC_5_133, I134=>output_MAC_5_134, I135=>output_MAC_5_135, I136=>output_MAC_5_136, I137=>output_MAC_5_137, I138=>output_MAC_5_138, I139=>output_MAC_5_139, I140=>output_MAC_5_140, I141=>output_MAC_5_141, I142=>output_MAC_5_142, I143=>output_MAC_5_143, I144=>output_MAC_5_144, I145=>output_MAC_5_145, I146=>output_MAC_5_146, I147=>output_MAC_5_147, I148=>output_MAC_5_148, I149=>output_MAC_5_149, I150=>output_MAC_5_150, I151=>output_MAC_5_151, I152=>output_MAC_5_152, I153=>output_MAC_5_153, I154=>output_MAC_5_154, I155=>output_MAC_5_155, I156=>output_MAC_5_156, I157=>output_MAC_5_157, I158=>output_MAC_5_158, I159=>output_MAC_5_159, I160=>output_MAC_5_160, I161=>output_MAC_5_161, I162=>output_MAC_5_162, I163=>output_MAC_5_163, I164=>output_MAC_5_164, I165=>output_MAC_5_165, I166=>output_MAC_5_166, I167=>output_MAC_5_167, I168=>output_MAC_5_168, I169=>output_MAC_5_169, I170=>output_MAC_5_170, I171=>output_MAC_5_171, I172=>output_MAC_5_172, I173=>output_MAC_5_173, I174=>output_MAC_5_174, I175=>output_MAC_5_175, I176=>output_MAC_5_176, I177=>output_MAC_5_177, I178=>output_MAC_5_178, I179=>output_MAC_5_179, I180=>output_MAC_5_180, I181=>output_MAC_5_181, I182=>output_MAC_5_182, I183=>output_MAC_5_183, I184=>output_MAC_5_184, I185=>output_MAC_5_185, I186=>output_MAC_5_186, I187=>output_MAC_5_187, I188=>output_MAC_5_188, I189=>output_MAC_5_189, I190=>output_MAC_5_190, I191=>output_MAC_5_191, I192=>output_MAC_5_192, I193=>output_MAC_5_193, I194=>output_MAC_5_194, I195=>output_MAC_5_195, I196=>output_MAC_5_196, I197=>output_MAC_5_197, I198=>output_MAC_5_198, I199=>output_MAC_5_199, I200=>output_MAC_5_200, I201=>output_MAC_5_201, I202=>output_MAC_5_202, I203=>output_MAC_5_203, I204=>output_MAC_5_204, I205=>output_MAC_5_205, I206=>output_MAC_5_206, I207=>output_MAC_5_207, I208=>output_MAC_5_208, I209=>output_MAC_5_209, I210=>output_MAC_5_210, I211=>output_MAC_5_211, I212=>output_MAC_5_212, I213=>output_MAC_5_213, I214=>output_MAC_5_214, I215=>output_MAC_5_215, I216=>output_MAC_5_216, I217=>output_MAC_5_217, I218=>output_MAC_5_218, I219=>output_MAC_5_219, I220=>output_MAC_5_220, I221=>output_MAC_5_221, I222=>output_MAC_5_222, I223=>output_MAC_5_223, I224=>output_MAC_5_224, I225=>output_MAC_5_225, I226=>output_MAC_5_226, I227=>output_MAC_5_227, I228=>output_MAC_5_228, I229=>output_MAC_5_229, I230=>output_MAC_5_230, I231=>output_MAC_5_231, I232=>output_MAC_5_232, I233=>output_MAC_5_233, I234=>output_MAC_5_234, I235=>output_MAC_5_235, I236=>output_MAC_5_236, I237=>output_MAC_5_237, I238=>output_MAC_5_238, I239=>output_MAC_5_239, I240=>output_MAC_5_240, I241=>output_MAC_5_241, I242=>output_MAC_5_242, I243=>output_MAC_5_243, I244=>output_MAC_5_244, I245=>output_MAC_5_245, I246=>output_MAC_5_246, I247=>output_MAC_5_247, I248=>output_MAC_5_248, I249=>output_MAC_5_249, I250=>output_MAC_5_250, I251=>output_MAC_5_251, I252=>output_MAC_5_252, I253=>output_MAC_5_253, I254=>output_MAC_5_254, I255=>output_MAC_5_255, I256=>output_MAC_5_256, I257=>output_MAC_5_257, I258=>output_MAC_5_258, I259=>output_MAC_5_259, I260=>output_MAC_5_260, I261=>output_MAC_5_261, I262=>output_MAC_5_262, I263=>output_MAC_5_263, I264=>output_MAC_5_264, I265=>output_MAC_5_265, I266=>output_MAC_5_266, I267=>output_MAC_5_267, I268=>output_MAC_5_268, I269=>output_MAC_5_269, I270=>output_MAC_5_270, I271=>output_MAC_5_271, I272=>output_MAC_5_272, I273=>output_MAC_5_273, I274=>output_MAC_5_274, I275=>output_MAC_5_275, I276=>output_MAC_5_276, I277=>output_MAC_5_277, I278=>output_MAC_5_278, I279=>output_MAC_5_279, I280=>output_MAC_5_280, I281=>output_MAC_5_281, I282=>output_MAC_5_282, I283=>output_MAC_5_283, I284=>output_MAC_5_284, I285=>output_MAC_5_285, I286=>output_MAC_5_286, I287=>output_MAC_5_287, I288=>output_MAC_5_288, I289=>output_MAC_5_289, I290=>output_MAC_5_290, I291=>output_MAC_5_291, I292=>output_MAC_5_292, I293=>output_MAC_5_293, I294=>output_MAC_5_294, I295=>output_MAC_5_295, I296=>output_MAC_5_296, I297=>output_MAC_5_297, I298=>output_MAC_5_298, I299=>output_MAC_5_299, I300=>output_MAC_5_300, I301=>output_MAC_5_301, I302=>output_MAC_5_302, I303=>output_MAC_5_303, I304=>output_MAC_5_304, I305=>output_MAC_5_305, I306=>output_MAC_5_306, I307=>output_MAC_5_307, I308=>output_MAC_5_308, I309=>output_MAC_5_309, I310=>output_MAC_5_310, I311=>output_MAC_5_311, I312=>output_MAC_5_312, I313=>output_MAC_5_313, I314=>output_MAC_5_314, I315=>output_MAC_5_315, I316=>output_MAC_5_316, I317=>output_MAC_5_317, I318=>output_MAC_5_318, I319=>output_MAC_5_319, I320=>output_MAC_5_320, I321=>output_MAC_5_321, I322=>output_MAC_5_322, I323=>output_MAC_5_323, I324=>output_MAC_5_324, I325=>output_MAC_5_325, I326=>output_MAC_5_326, I327=>output_MAC_5_327, I328=>output_MAC_5_328, I329=>output_MAC_5_329, I330=>output_MAC_5_330, I331=>output_MAC_5_331, I332=>output_MAC_5_332, I333=>output_MAC_5_333, I334=>output_MAC_5_334, I335=>output_MAC_5_335, I336=>output_MAC_5_336, I337=>output_MAC_5_337, I338=>output_MAC_5_338, I339=>output_MAC_5_339, I340=>output_MAC_5_340, I341=>output_MAC_5_341, I342=>output_MAC_5_342, I343=>output_MAC_5_343, I344=>output_MAC_5_344, I345=>output_MAC_5_345, I346=>output_MAC_5_346, I347=>output_MAC_5_347, I348=>output_MAC_5_348, I349=>output_MAC_5_349, I350=>output_MAC_5_350, I351=>output_MAC_5_351, I352=>output_MAC_5_352, I353=>output_MAC_5_353, I354=>output_MAC_5_354, I355=>output_MAC_5_355, I356=>output_MAC_5_356, I357=>output_MAC_5_357, I358=>output_MAC_5_358, I359=>output_MAC_5_359, I360=>output_MAC_5_360, I361=>output_MAC_5_361, I362=>output_MAC_5_362, I363=>output_MAC_5_363, I364=>output_MAC_5_364, I365=>output_MAC_5_365, I366=>output_MAC_5_366, I367=>output_MAC_5_367, I368=>output_MAC_5_368, I369=>output_MAC_5_369, I370=>output_MAC_5_370, I371=>output_MAC_5_371, I372=>output_MAC_5_372, I373=>output_MAC_5_373, I374=>output_MAC_5_374, I375=>output_MAC_5_375, I376=>output_MAC_5_376, I377=>output_MAC_5_377, I378=>output_MAC_5_378, I379=>output_MAC_5_379, I380=>output_MAC_5_380, I381=>output_MAC_5_381, I382=>output_MAC_5_382, I383=>output_MAC_5_383, I384=>output_MAC_5_384, I385=>output_MAC_5_385, I386=>output_MAC_5_386, I387=>output_MAC_5_387, I388=>output_MAC_5_388, I389=>output_MAC_5_389, I390=>output_MAC_5_390, I391=>output_MAC_5_391, I392=>output_MAC_5_392, I393=>output_MAC_5_393, I394=>output_MAC_5_394, I395=>output_MAC_5_395, I396=>output_MAC_5_396, I397=>output_MAC_5_397, I398=>output_MAC_5_398, I399=>output_MAC_5_399, I400=>output_MAC_5_400, I401=>output_MAC_5_401, I402=>output_MAC_5_402, I403=>output_MAC_5_403, I404=>output_MAC_5_404, I405=>output_MAC_5_405, I406=>output_MAC_5_406, I407=>output_MAC_5_407, I408=>output_MAC_5_408, I409=>output_MAC_5_409, I410=>output_MAC_5_410, I411=>output_MAC_5_411, I412=>output_MAC_5_412, I413=>output_MAC_5_413, I414=>output_MAC_5_414, I415=>output_MAC_5_415, I416=>output_MAC_5_416, I417=>output_MAC_5_417, I418=>output_MAC_5_418, I419=>output_MAC_5_419, I420=>output_MAC_5_420, I421=>output_MAC_5_421, I422=>output_MAC_5_422, I423=>output_MAC_5_423, I424=>output_MAC_5_424, I425=>output_MAC_5_425, I426=>output_MAC_5_426, I427=>output_MAC_5_427, I428=>output_MAC_5_428, I429=>output_MAC_5_429, I430=>output_MAC_5_430, I431=>output_MAC_5_431, I432=>output_MAC_5_432, I433=>output_MAC_5_433, I434=>output_MAC_5_434, I435=>output_MAC_5_435, I436=>output_MAC_5_436, I437=>output_MAC_5_437, I438=>output_MAC_5_438, I439=>output_MAC_5_439, I440=>output_MAC_5_440, I441=>output_MAC_5_441, I442=>output_MAC_5_442, I443=>output_MAC_5_443, I444=>output_MAC_5_444, I445=>output_MAC_5_445, I446=>output_MAC_5_446, I447=>output_MAC_5_447, I448=>output_MAC_5_448, I449=>output_MAC_5_449, I450=>output_MAC_5_450, I451=>output_MAC_5_451, I452=>output_MAC_5_452, I453=>output_MAC_5_453, I454=>output_MAC_5_454, I455=>output_MAC_5_455, I456=>output_MAC_5_456, I457=>output_MAC_5_457, I458=>output_MAC_5_458, I459=>output_MAC_5_459, I460=>output_MAC_5_460, I461=>output_MAC_5_461, I462=>output_MAC_5_462, I463=>output_MAC_5_463, I464=>output_MAC_5_464, I465=>output_MAC_5_465, I466=>output_MAC_5_466, I467=>output_MAC_5_467, I468=>output_MAC_5_468, I469=>output_MAC_5_469, I470=>output_MAC_5_470, I471=>output_MAC_5_471, I472=>output_MAC_5_472, I473=>output_MAC_5_473, I474=>output_MAC_5_474, I475=>output_MAC_5_475, I476=>output_MAC_5_476, I477=>output_MAC_5_477, I478=>output_MAC_5_478, I479=>output_MAC_5_479, I480=>output_MAC_5_480, I481=>output_MAC_5_481, I482=>output_MAC_5_482, I483=>output_MAC_5_483, I484=>output_MAC_5_484, I485=>output_MAC_5_485, I486=>output_MAC_5_486, I487=>output_MAC_5_487, I488=>output_MAC_5_488, I489=>output_MAC_5_489, I490=>output_MAC_5_490, I491=>output_MAC_5_491, I492=>output_MAC_5_492, I493=>output_MAC_5_493, I494=>output_MAC_5_494, I495=>output_MAC_5_495, I496=>output_MAC_5_496, I497=>output_MAC_5_497, I498=>output_MAC_5_498, I499=>output_MAC_5_499, I500=>output_MAC_5_500, I501=>output_MAC_5_501, I502=>output_MAC_5_502, I503=>output_MAC_5_503, I504=>output_MAC_5_504, I505=>output_MAC_5_505, I506=>output_MAC_5_506, I507=>output_MAC_5_507, I508=>output_MAC_5_508, I509=>output_MAC_5_509, I510=>output_MAC_5_510, I511=>output_MAC_5_511, I512=>output_MAC_5_512, I513=>output_MAC_5_513, I514=>output_MAC_5_514, I515=>output_MAC_5_515, I516=>output_MAC_5_516, I517=>output_MAC_5_517, I518=>output_MAC_5_518, I519=>output_MAC_5_519, I520=>output_MAC_5_520, I521=>output_MAC_5_521, I522=>output_MAC_5_522, I523=>output_MAC_5_523, I524=>output_MAC_5_524, I525=>output_MAC_5_525, I526=>output_MAC_5_526, I527=>output_MAC_5_527, I528=>output_MAC_5_528, I529=>output_MAC_5_529, I530=>output_MAC_5_530, I531=>output_MAC_5_531, I532=>output_MAC_5_532, I533=>output_MAC_5_533, I534=>output_MAC_5_534, I535=>output_MAC_5_535, I536=>output_MAC_5_536, I537=>output_MAC_5_537, I538=>output_MAC_5_538, I539=>output_MAC_5_539, I540=>output_MAC_5_540, I541=>output_MAC_5_541, I542=>output_MAC_5_542, I543=>output_MAC_5_543, I544=>output_MAC_5_544, I545=>output_MAC_5_545, I546=>output_MAC_5_546, I547=>output_MAC_5_547, I548=>output_MAC_5_548, I549=>output_MAC_5_549, I550=>output_MAC_5_550, I551=>output_MAC_5_551, I552=>output_MAC_5_552, I553=>output_MAC_5_553, I554=>output_MAC_5_554, I555=>output_MAC_5_555, I556=>output_MAC_5_556, I557=>output_MAC_5_557, I558=>output_MAC_5_558, I559=>output_MAC_5_559, I560=>output_MAC_5_560, I561=>output_MAC_5_561, I562=>output_MAC_5_562, I563=>output_MAC_5_563, I564=>output_MAC_5_564, I565=>output_MAC_5_565, I566=>output_MAC_5_566, I567=>output_MAC_5_567, I568=>output_MAC_5_568, I569=>output_MAC_5_569, I570=>output_MAC_5_570, I571=>output_MAC_5_571, I572=>output_MAC_5_572, I573=>output_MAC_5_573, I574=>output_MAC_5_574, I575=>output_MAC_5_575, I576=>output_MAC_5_576, I577=>output_MAC_5_577, I578=>output_MAC_5_578, I579=>output_MAC_5_579, I580=>output_MAC_5_580, I581=>output_MAC_5_581, I582=>output_MAC_5_582, I583=>output_MAC_5_583, I584=>output_MAC_5_584, I585=>output_MAC_5_585, I586=>output_MAC_5_586, I587=>output_MAC_5_587, I588=>output_MAC_5_588, I589=>output_MAC_5_589, I590=>output_MAC_5_590, I591=>output_MAC_5_591, I592=>output_MAC_5_592, I593=>output_MAC_5_593, I594=>output_MAC_5_594, I595=>output_MAC_5_595, I596=>output_MAC_5_596, I597=>output_MAC_5_597, I598=>output_MAC_5_598, I599=>output_MAC_5_599, I600=>output_MAC_5_600, I601=>output_MAC_5_601, I602=>output_MAC_5_602, I603=>output_MAC_5_603, I604=>output_MAC_5_604, I605=>output_MAC_5_605, I606=>output_MAC_5_606, I607=>output_MAC_5_607, I608=>output_MAC_5_608, I609=>output_MAC_5_609, I610=>output_MAC_5_610, I611=>output_MAC_5_611, I612=>output_MAC_5_612, I613=>output_MAC_5_613, I614=>output_MAC_5_614, I615=>output_MAC_5_615, I616=>output_MAC_5_616, I617=>output_MAC_5_617, I618=>output_MAC_5_618, I619=>output_MAC_5_619, I620=>output_MAC_5_620, I621=>output_MAC_5_621, I622=>output_MAC_5_622, I623=>output_MAC_5_623, I624=>output_MAC_5_624, I625=>output_MAC_5_625, I626=>output_MAC_5_626, I627=>output_MAC_5_627, I628=>output_MAC_5_628, I629=>output_MAC_5_629, I630=>output_MAC_5_630, I631=>output_MAC_5_631, I632=>output_MAC_5_632, I633=>output_MAC_5_633, I634=>output_MAC_5_634, I635=>output_MAC_5_635, I636=>output_MAC_5_636, I637=>output_MAC_5_637, I638=>output_MAC_5_638, I639=>output_MAC_5_639, I640=>output_MAC_5_640, I641=>output_MAC_5_641, I642=>output_MAC_5_642, I643=>output_MAC_5_643, I644=>output_MAC_5_644, I645=>output_MAC_5_645, I646=>output_MAC_5_646, I647=>output_MAC_5_647, I648=>output_MAC_5_648, I649=>output_MAC_5_649, I650=>output_MAC_5_650, I651=>output_MAC_5_651, I652=>output_MAC_5_652, I653=>output_MAC_5_653, I654=>output_MAC_5_654, I655=>output_MAC_5_655, I656=>output_MAC_5_656, I657=>output_MAC_5_657, I658=>output_MAC_5_658, I659=>output_MAC_5_659, I660=>output_MAC_5_660, I661=>output_MAC_5_661, I662=>output_MAC_5_662, I663=>output_MAC_5_663, I664=>output_MAC_5_664, I665=>output_MAC_5_665, I666=>output_MAC_5_666, I667=>output_MAC_5_667, I668=>output_MAC_5_668, I669=>output_MAC_5_669, I670=>output_MAC_5_670, I671=>output_MAC_5_671, I672=>output_MAC_5_672, I673=>output_MAC_5_673, I674=>output_MAC_5_674, I675=>output_MAC_5_675, I676=>output_MAC_5_676, I677=>output_MAC_5_677, I678=>output_MAC_5_678, I679=>output_MAC_5_679, I680=>output_MAC_5_680, I681=>output_MAC_5_681, I682=>output_MAC_5_682, I683=>output_MAC_5_683, I684=>output_MAC_5_684, I685=>output_MAC_5_685, I686=>output_MAC_5_686, I687=>output_MAC_5_687, I688=>output_MAC_5_688, I689=>output_MAC_5_689, I690=>output_MAC_5_690, I691=>output_MAC_5_691, I692=>output_MAC_5_692, I693=>output_MAC_5_693, I694=>output_MAC_5_694, I695=>output_MAC_5_695, I696=>output_MAC_5_696, I697=>output_MAC_5_697, I698=>output_MAC_5_698, I699=>output_MAC_5_699, I700=>output_MAC_5_700, I701=>output_MAC_5_701, I702=>output_MAC_5_702, I703=>output_MAC_5_703, I704=>output_MAC_5_704, I705=>output_MAC_5_705, I706=>output_MAC_5_706, I707=>output_MAC_5_707, I708=>output_MAC_5_708, I709=>output_MAC_5_709, I710=>output_MAC_5_710, I711=>output_MAC_5_711, I712=>output_MAC_5_712, I713=>output_MAC_5_713, I714=>output_MAC_5_714, I715=>output_MAC_5_715, I716=>output_MAC_5_716, I717=>output_MAC_5_717, I718=>output_MAC_5_718, I719=>output_MAC_5_719, I720=>output_MAC_5_720, I721=>output_MAC_5_721, I722=>output_MAC_5_722, I723=>output_MAC_5_723, I724=>output_MAC_5_724, I725=>output_MAC_5_725, I726=>output_MAC_5_726, I727=>output_MAC_5_727, I728=>output_MAC_5_728, I729=>output_MAC_5_729, I730=>output_MAC_5_730, I731=>output_MAC_5_731, I732=>output_MAC_5_732, I733=>output_MAC_5_733, I734=>output_MAC_5_734, I735=>output_MAC_5_735, I736=>output_MAC_5_736, I737=>output_MAC_5_737, I738=>output_MAC_5_738, I739=>output_MAC_5_739, I740=>output_MAC_5_740, I741=>output_MAC_5_741, I742=>output_MAC_5_742, I743=>output_MAC_5_743, I744=>output_MAC_5_744, I745=>output_MAC_5_745, I746=>output_MAC_5_746, I747=>output_MAC_5_747, I748=>output_MAC_5_748, I749=>output_MAC_5_749, I750=>output_MAC_5_750, I751=>output_MAC_5_751, I752=>output_MAC_5_752, I753=>output_MAC_5_753, I754=>output_MAC_5_754, I755=>output_MAC_5_755, I756=>output_MAC_5_756, I757=>output_MAC_5_757, I758=>output_MAC_5_758, I759=>output_MAC_5_759, I760=>output_MAC_5_760, I761=>output_MAC_5_761, I762=>output_MAC_5_762, I763=>output_MAC_5_763, I764=>output_MAC_5_764, I765=>output_MAC_5_765, I766=>output_MAC_5_766, I767=>output_MAC_5_767, 
		SEL_mux=>SEL_mux, O=>output_row_5);

	mux_row_6: mux_768to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_6_0, I1=>output_MAC_6_1, I2=>output_MAC_6_2, I3=>output_MAC_6_3, I4=>output_MAC_6_4, I5=>output_MAC_6_5, I6=>output_MAC_6_6, I7=>output_MAC_6_7, I8=>output_MAC_6_8, I9=>output_MAC_6_9, I10=>output_MAC_6_10, I11=>output_MAC_6_11, I12=>output_MAC_6_12, I13=>output_MAC_6_13, I14=>output_MAC_6_14, I15=>output_MAC_6_15, I16=>output_MAC_6_16, I17=>output_MAC_6_17, I18=>output_MAC_6_18, I19=>output_MAC_6_19, I20=>output_MAC_6_20, I21=>output_MAC_6_21, I22=>output_MAC_6_22, I23=>output_MAC_6_23, I24=>output_MAC_6_24, I25=>output_MAC_6_25, I26=>output_MAC_6_26, I27=>output_MAC_6_27, I28=>output_MAC_6_28, I29=>output_MAC_6_29, I30=>output_MAC_6_30, I31=>output_MAC_6_31, I32=>output_MAC_6_32, I33=>output_MAC_6_33, I34=>output_MAC_6_34, I35=>output_MAC_6_35, I36=>output_MAC_6_36, I37=>output_MAC_6_37, I38=>output_MAC_6_38, I39=>output_MAC_6_39, I40=>output_MAC_6_40, I41=>output_MAC_6_41, I42=>output_MAC_6_42, I43=>output_MAC_6_43, I44=>output_MAC_6_44, I45=>output_MAC_6_45, I46=>output_MAC_6_46, I47=>output_MAC_6_47, I48=>output_MAC_6_48, I49=>output_MAC_6_49, I50=>output_MAC_6_50, I51=>output_MAC_6_51, I52=>output_MAC_6_52, I53=>output_MAC_6_53, I54=>output_MAC_6_54, I55=>output_MAC_6_55, I56=>output_MAC_6_56, I57=>output_MAC_6_57, I58=>output_MAC_6_58, I59=>output_MAC_6_59, I60=>output_MAC_6_60, I61=>output_MAC_6_61, I62=>output_MAC_6_62, I63=>output_MAC_6_63, I64=>output_MAC_6_64, I65=>output_MAC_6_65, I66=>output_MAC_6_66, I67=>output_MAC_6_67, I68=>output_MAC_6_68, I69=>output_MAC_6_69, I70=>output_MAC_6_70, I71=>output_MAC_6_71, I72=>output_MAC_6_72, I73=>output_MAC_6_73, I74=>output_MAC_6_74, I75=>output_MAC_6_75, I76=>output_MAC_6_76, I77=>output_MAC_6_77, I78=>output_MAC_6_78, I79=>output_MAC_6_79, I80=>output_MAC_6_80, I81=>output_MAC_6_81, I82=>output_MAC_6_82, I83=>output_MAC_6_83, I84=>output_MAC_6_84, I85=>output_MAC_6_85, I86=>output_MAC_6_86, I87=>output_MAC_6_87, I88=>output_MAC_6_88, I89=>output_MAC_6_89, I90=>output_MAC_6_90, I91=>output_MAC_6_91, I92=>output_MAC_6_92, I93=>output_MAC_6_93, I94=>output_MAC_6_94, I95=>output_MAC_6_95, I96=>output_MAC_6_96, I97=>output_MAC_6_97, I98=>output_MAC_6_98, I99=>output_MAC_6_99, I100=>output_MAC_6_100, I101=>output_MAC_6_101, I102=>output_MAC_6_102, I103=>output_MAC_6_103, I104=>output_MAC_6_104, I105=>output_MAC_6_105, I106=>output_MAC_6_106, I107=>output_MAC_6_107, I108=>output_MAC_6_108, I109=>output_MAC_6_109, I110=>output_MAC_6_110, I111=>output_MAC_6_111, I112=>output_MAC_6_112, I113=>output_MAC_6_113, I114=>output_MAC_6_114, I115=>output_MAC_6_115, I116=>output_MAC_6_116, I117=>output_MAC_6_117, I118=>output_MAC_6_118, I119=>output_MAC_6_119, I120=>output_MAC_6_120, I121=>output_MAC_6_121, I122=>output_MAC_6_122, I123=>output_MAC_6_123, I124=>output_MAC_6_124, I125=>output_MAC_6_125, I126=>output_MAC_6_126, I127=>output_MAC_6_127, I128=>output_MAC_6_128, I129=>output_MAC_6_129, I130=>output_MAC_6_130, I131=>output_MAC_6_131, I132=>output_MAC_6_132, I133=>output_MAC_6_133, I134=>output_MAC_6_134, I135=>output_MAC_6_135, I136=>output_MAC_6_136, I137=>output_MAC_6_137, I138=>output_MAC_6_138, I139=>output_MAC_6_139, I140=>output_MAC_6_140, I141=>output_MAC_6_141, I142=>output_MAC_6_142, I143=>output_MAC_6_143, I144=>output_MAC_6_144, I145=>output_MAC_6_145, I146=>output_MAC_6_146, I147=>output_MAC_6_147, I148=>output_MAC_6_148, I149=>output_MAC_6_149, I150=>output_MAC_6_150, I151=>output_MAC_6_151, I152=>output_MAC_6_152, I153=>output_MAC_6_153, I154=>output_MAC_6_154, I155=>output_MAC_6_155, I156=>output_MAC_6_156, I157=>output_MAC_6_157, I158=>output_MAC_6_158, I159=>output_MAC_6_159, I160=>output_MAC_6_160, I161=>output_MAC_6_161, I162=>output_MAC_6_162, I163=>output_MAC_6_163, I164=>output_MAC_6_164, I165=>output_MAC_6_165, I166=>output_MAC_6_166, I167=>output_MAC_6_167, I168=>output_MAC_6_168, I169=>output_MAC_6_169, I170=>output_MAC_6_170, I171=>output_MAC_6_171, I172=>output_MAC_6_172, I173=>output_MAC_6_173, I174=>output_MAC_6_174, I175=>output_MAC_6_175, I176=>output_MAC_6_176, I177=>output_MAC_6_177, I178=>output_MAC_6_178, I179=>output_MAC_6_179, I180=>output_MAC_6_180, I181=>output_MAC_6_181, I182=>output_MAC_6_182, I183=>output_MAC_6_183, I184=>output_MAC_6_184, I185=>output_MAC_6_185, I186=>output_MAC_6_186, I187=>output_MAC_6_187, I188=>output_MAC_6_188, I189=>output_MAC_6_189, I190=>output_MAC_6_190, I191=>output_MAC_6_191, I192=>output_MAC_6_192, I193=>output_MAC_6_193, I194=>output_MAC_6_194, I195=>output_MAC_6_195, I196=>output_MAC_6_196, I197=>output_MAC_6_197, I198=>output_MAC_6_198, I199=>output_MAC_6_199, I200=>output_MAC_6_200, I201=>output_MAC_6_201, I202=>output_MAC_6_202, I203=>output_MAC_6_203, I204=>output_MAC_6_204, I205=>output_MAC_6_205, I206=>output_MAC_6_206, I207=>output_MAC_6_207, I208=>output_MAC_6_208, I209=>output_MAC_6_209, I210=>output_MAC_6_210, I211=>output_MAC_6_211, I212=>output_MAC_6_212, I213=>output_MAC_6_213, I214=>output_MAC_6_214, I215=>output_MAC_6_215, I216=>output_MAC_6_216, I217=>output_MAC_6_217, I218=>output_MAC_6_218, I219=>output_MAC_6_219, I220=>output_MAC_6_220, I221=>output_MAC_6_221, I222=>output_MAC_6_222, I223=>output_MAC_6_223, I224=>output_MAC_6_224, I225=>output_MAC_6_225, I226=>output_MAC_6_226, I227=>output_MAC_6_227, I228=>output_MAC_6_228, I229=>output_MAC_6_229, I230=>output_MAC_6_230, I231=>output_MAC_6_231, I232=>output_MAC_6_232, I233=>output_MAC_6_233, I234=>output_MAC_6_234, I235=>output_MAC_6_235, I236=>output_MAC_6_236, I237=>output_MAC_6_237, I238=>output_MAC_6_238, I239=>output_MAC_6_239, I240=>output_MAC_6_240, I241=>output_MAC_6_241, I242=>output_MAC_6_242, I243=>output_MAC_6_243, I244=>output_MAC_6_244, I245=>output_MAC_6_245, I246=>output_MAC_6_246, I247=>output_MAC_6_247, I248=>output_MAC_6_248, I249=>output_MAC_6_249, I250=>output_MAC_6_250, I251=>output_MAC_6_251, I252=>output_MAC_6_252, I253=>output_MAC_6_253, I254=>output_MAC_6_254, I255=>output_MAC_6_255, I256=>output_MAC_6_256, I257=>output_MAC_6_257, I258=>output_MAC_6_258, I259=>output_MAC_6_259, I260=>output_MAC_6_260, I261=>output_MAC_6_261, I262=>output_MAC_6_262, I263=>output_MAC_6_263, I264=>output_MAC_6_264, I265=>output_MAC_6_265, I266=>output_MAC_6_266, I267=>output_MAC_6_267, I268=>output_MAC_6_268, I269=>output_MAC_6_269, I270=>output_MAC_6_270, I271=>output_MAC_6_271, I272=>output_MAC_6_272, I273=>output_MAC_6_273, I274=>output_MAC_6_274, I275=>output_MAC_6_275, I276=>output_MAC_6_276, I277=>output_MAC_6_277, I278=>output_MAC_6_278, I279=>output_MAC_6_279, I280=>output_MAC_6_280, I281=>output_MAC_6_281, I282=>output_MAC_6_282, I283=>output_MAC_6_283, I284=>output_MAC_6_284, I285=>output_MAC_6_285, I286=>output_MAC_6_286, I287=>output_MAC_6_287, I288=>output_MAC_6_288, I289=>output_MAC_6_289, I290=>output_MAC_6_290, I291=>output_MAC_6_291, I292=>output_MAC_6_292, I293=>output_MAC_6_293, I294=>output_MAC_6_294, I295=>output_MAC_6_295, I296=>output_MAC_6_296, I297=>output_MAC_6_297, I298=>output_MAC_6_298, I299=>output_MAC_6_299, I300=>output_MAC_6_300, I301=>output_MAC_6_301, I302=>output_MAC_6_302, I303=>output_MAC_6_303, I304=>output_MAC_6_304, I305=>output_MAC_6_305, I306=>output_MAC_6_306, I307=>output_MAC_6_307, I308=>output_MAC_6_308, I309=>output_MAC_6_309, I310=>output_MAC_6_310, I311=>output_MAC_6_311, I312=>output_MAC_6_312, I313=>output_MAC_6_313, I314=>output_MAC_6_314, I315=>output_MAC_6_315, I316=>output_MAC_6_316, I317=>output_MAC_6_317, I318=>output_MAC_6_318, I319=>output_MAC_6_319, I320=>output_MAC_6_320, I321=>output_MAC_6_321, I322=>output_MAC_6_322, I323=>output_MAC_6_323, I324=>output_MAC_6_324, I325=>output_MAC_6_325, I326=>output_MAC_6_326, I327=>output_MAC_6_327, I328=>output_MAC_6_328, I329=>output_MAC_6_329, I330=>output_MAC_6_330, I331=>output_MAC_6_331, I332=>output_MAC_6_332, I333=>output_MAC_6_333, I334=>output_MAC_6_334, I335=>output_MAC_6_335, I336=>output_MAC_6_336, I337=>output_MAC_6_337, I338=>output_MAC_6_338, I339=>output_MAC_6_339, I340=>output_MAC_6_340, I341=>output_MAC_6_341, I342=>output_MAC_6_342, I343=>output_MAC_6_343, I344=>output_MAC_6_344, I345=>output_MAC_6_345, I346=>output_MAC_6_346, I347=>output_MAC_6_347, I348=>output_MAC_6_348, I349=>output_MAC_6_349, I350=>output_MAC_6_350, I351=>output_MAC_6_351, I352=>output_MAC_6_352, I353=>output_MAC_6_353, I354=>output_MAC_6_354, I355=>output_MAC_6_355, I356=>output_MAC_6_356, I357=>output_MAC_6_357, I358=>output_MAC_6_358, I359=>output_MAC_6_359, I360=>output_MAC_6_360, I361=>output_MAC_6_361, I362=>output_MAC_6_362, I363=>output_MAC_6_363, I364=>output_MAC_6_364, I365=>output_MAC_6_365, I366=>output_MAC_6_366, I367=>output_MAC_6_367, I368=>output_MAC_6_368, I369=>output_MAC_6_369, I370=>output_MAC_6_370, I371=>output_MAC_6_371, I372=>output_MAC_6_372, I373=>output_MAC_6_373, I374=>output_MAC_6_374, I375=>output_MAC_6_375, I376=>output_MAC_6_376, I377=>output_MAC_6_377, I378=>output_MAC_6_378, I379=>output_MAC_6_379, I380=>output_MAC_6_380, I381=>output_MAC_6_381, I382=>output_MAC_6_382, I383=>output_MAC_6_383, I384=>output_MAC_6_384, I385=>output_MAC_6_385, I386=>output_MAC_6_386, I387=>output_MAC_6_387, I388=>output_MAC_6_388, I389=>output_MAC_6_389, I390=>output_MAC_6_390, I391=>output_MAC_6_391, I392=>output_MAC_6_392, I393=>output_MAC_6_393, I394=>output_MAC_6_394, I395=>output_MAC_6_395, I396=>output_MAC_6_396, I397=>output_MAC_6_397, I398=>output_MAC_6_398, I399=>output_MAC_6_399, I400=>output_MAC_6_400, I401=>output_MAC_6_401, I402=>output_MAC_6_402, I403=>output_MAC_6_403, I404=>output_MAC_6_404, I405=>output_MAC_6_405, I406=>output_MAC_6_406, I407=>output_MAC_6_407, I408=>output_MAC_6_408, I409=>output_MAC_6_409, I410=>output_MAC_6_410, I411=>output_MAC_6_411, I412=>output_MAC_6_412, I413=>output_MAC_6_413, I414=>output_MAC_6_414, I415=>output_MAC_6_415, I416=>output_MAC_6_416, I417=>output_MAC_6_417, I418=>output_MAC_6_418, I419=>output_MAC_6_419, I420=>output_MAC_6_420, I421=>output_MAC_6_421, I422=>output_MAC_6_422, I423=>output_MAC_6_423, I424=>output_MAC_6_424, I425=>output_MAC_6_425, I426=>output_MAC_6_426, I427=>output_MAC_6_427, I428=>output_MAC_6_428, I429=>output_MAC_6_429, I430=>output_MAC_6_430, I431=>output_MAC_6_431, I432=>output_MAC_6_432, I433=>output_MAC_6_433, I434=>output_MAC_6_434, I435=>output_MAC_6_435, I436=>output_MAC_6_436, I437=>output_MAC_6_437, I438=>output_MAC_6_438, I439=>output_MAC_6_439, I440=>output_MAC_6_440, I441=>output_MAC_6_441, I442=>output_MAC_6_442, I443=>output_MAC_6_443, I444=>output_MAC_6_444, I445=>output_MAC_6_445, I446=>output_MAC_6_446, I447=>output_MAC_6_447, I448=>output_MAC_6_448, I449=>output_MAC_6_449, I450=>output_MAC_6_450, I451=>output_MAC_6_451, I452=>output_MAC_6_452, I453=>output_MAC_6_453, I454=>output_MAC_6_454, I455=>output_MAC_6_455, I456=>output_MAC_6_456, I457=>output_MAC_6_457, I458=>output_MAC_6_458, I459=>output_MAC_6_459, I460=>output_MAC_6_460, I461=>output_MAC_6_461, I462=>output_MAC_6_462, I463=>output_MAC_6_463, I464=>output_MAC_6_464, I465=>output_MAC_6_465, I466=>output_MAC_6_466, I467=>output_MAC_6_467, I468=>output_MAC_6_468, I469=>output_MAC_6_469, I470=>output_MAC_6_470, I471=>output_MAC_6_471, I472=>output_MAC_6_472, I473=>output_MAC_6_473, I474=>output_MAC_6_474, I475=>output_MAC_6_475, I476=>output_MAC_6_476, I477=>output_MAC_6_477, I478=>output_MAC_6_478, I479=>output_MAC_6_479, I480=>output_MAC_6_480, I481=>output_MAC_6_481, I482=>output_MAC_6_482, I483=>output_MAC_6_483, I484=>output_MAC_6_484, I485=>output_MAC_6_485, I486=>output_MAC_6_486, I487=>output_MAC_6_487, I488=>output_MAC_6_488, I489=>output_MAC_6_489, I490=>output_MAC_6_490, I491=>output_MAC_6_491, I492=>output_MAC_6_492, I493=>output_MAC_6_493, I494=>output_MAC_6_494, I495=>output_MAC_6_495, I496=>output_MAC_6_496, I497=>output_MAC_6_497, I498=>output_MAC_6_498, I499=>output_MAC_6_499, I500=>output_MAC_6_500, I501=>output_MAC_6_501, I502=>output_MAC_6_502, I503=>output_MAC_6_503, I504=>output_MAC_6_504, I505=>output_MAC_6_505, I506=>output_MAC_6_506, I507=>output_MAC_6_507, I508=>output_MAC_6_508, I509=>output_MAC_6_509, I510=>output_MAC_6_510, I511=>output_MAC_6_511, I512=>output_MAC_6_512, I513=>output_MAC_6_513, I514=>output_MAC_6_514, I515=>output_MAC_6_515, I516=>output_MAC_6_516, I517=>output_MAC_6_517, I518=>output_MAC_6_518, I519=>output_MAC_6_519, I520=>output_MAC_6_520, I521=>output_MAC_6_521, I522=>output_MAC_6_522, I523=>output_MAC_6_523, I524=>output_MAC_6_524, I525=>output_MAC_6_525, I526=>output_MAC_6_526, I527=>output_MAC_6_527, I528=>output_MAC_6_528, I529=>output_MAC_6_529, I530=>output_MAC_6_530, I531=>output_MAC_6_531, I532=>output_MAC_6_532, I533=>output_MAC_6_533, I534=>output_MAC_6_534, I535=>output_MAC_6_535, I536=>output_MAC_6_536, I537=>output_MAC_6_537, I538=>output_MAC_6_538, I539=>output_MAC_6_539, I540=>output_MAC_6_540, I541=>output_MAC_6_541, I542=>output_MAC_6_542, I543=>output_MAC_6_543, I544=>output_MAC_6_544, I545=>output_MAC_6_545, I546=>output_MAC_6_546, I547=>output_MAC_6_547, I548=>output_MAC_6_548, I549=>output_MAC_6_549, I550=>output_MAC_6_550, I551=>output_MAC_6_551, I552=>output_MAC_6_552, I553=>output_MAC_6_553, I554=>output_MAC_6_554, I555=>output_MAC_6_555, I556=>output_MAC_6_556, I557=>output_MAC_6_557, I558=>output_MAC_6_558, I559=>output_MAC_6_559, I560=>output_MAC_6_560, I561=>output_MAC_6_561, I562=>output_MAC_6_562, I563=>output_MAC_6_563, I564=>output_MAC_6_564, I565=>output_MAC_6_565, I566=>output_MAC_6_566, I567=>output_MAC_6_567, I568=>output_MAC_6_568, I569=>output_MAC_6_569, I570=>output_MAC_6_570, I571=>output_MAC_6_571, I572=>output_MAC_6_572, I573=>output_MAC_6_573, I574=>output_MAC_6_574, I575=>output_MAC_6_575, I576=>output_MAC_6_576, I577=>output_MAC_6_577, I578=>output_MAC_6_578, I579=>output_MAC_6_579, I580=>output_MAC_6_580, I581=>output_MAC_6_581, I582=>output_MAC_6_582, I583=>output_MAC_6_583, I584=>output_MAC_6_584, I585=>output_MAC_6_585, I586=>output_MAC_6_586, I587=>output_MAC_6_587, I588=>output_MAC_6_588, I589=>output_MAC_6_589, I590=>output_MAC_6_590, I591=>output_MAC_6_591, I592=>output_MAC_6_592, I593=>output_MAC_6_593, I594=>output_MAC_6_594, I595=>output_MAC_6_595, I596=>output_MAC_6_596, I597=>output_MAC_6_597, I598=>output_MAC_6_598, I599=>output_MAC_6_599, I600=>output_MAC_6_600, I601=>output_MAC_6_601, I602=>output_MAC_6_602, I603=>output_MAC_6_603, I604=>output_MAC_6_604, I605=>output_MAC_6_605, I606=>output_MAC_6_606, I607=>output_MAC_6_607, I608=>output_MAC_6_608, I609=>output_MAC_6_609, I610=>output_MAC_6_610, I611=>output_MAC_6_611, I612=>output_MAC_6_612, I613=>output_MAC_6_613, I614=>output_MAC_6_614, I615=>output_MAC_6_615, I616=>output_MAC_6_616, I617=>output_MAC_6_617, I618=>output_MAC_6_618, I619=>output_MAC_6_619, I620=>output_MAC_6_620, I621=>output_MAC_6_621, I622=>output_MAC_6_622, I623=>output_MAC_6_623, I624=>output_MAC_6_624, I625=>output_MAC_6_625, I626=>output_MAC_6_626, I627=>output_MAC_6_627, I628=>output_MAC_6_628, I629=>output_MAC_6_629, I630=>output_MAC_6_630, I631=>output_MAC_6_631, I632=>output_MAC_6_632, I633=>output_MAC_6_633, I634=>output_MAC_6_634, I635=>output_MAC_6_635, I636=>output_MAC_6_636, I637=>output_MAC_6_637, I638=>output_MAC_6_638, I639=>output_MAC_6_639, I640=>output_MAC_6_640, I641=>output_MAC_6_641, I642=>output_MAC_6_642, I643=>output_MAC_6_643, I644=>output_MAC_6_644, I645=>output_MAC_6_645, I646=>output_MAC_6_646, I647=>output_MAC_6_647, I648=>output_MAC_6_648, I649=>output_MAC_6_649, I650=>output_MAC_6_650, I651=>output_MAC_6_651, I652=>output_MAC_6_652, I653=>output_MAC_6_653, I654=>output_MAC_6_654, I655=>output_MAC_6_655, I656=>output_MAC_6_656, I657=>output_MAC_6_657, I658=>output_MAC_6_658, I659=>output_MAC_6_659, I660=>output_MAC_6_660, I661=>output_MAC_6_661, I662=>output_MAC_6_662, I663=>output_MAC_6_663, I664=>output_MAC_6_664, I665=>output_MAC_6_665, I666=>output_MAC_6_666, I667=>output_MAC_6_667, I668=>output_MAC_6_668, I669=>output_MAC_6_669, I670=>output_MAC_6_670, I671=>output_MAC_6_671, I672=>output_MAC_6_672, I673=>output_MAC_6_673, I674=>output_MAC_6_674, I675=>output_MAC_6_675, I676=>output_MAC_6_676, I677=>output_MAC_6_677, I678=>output_MAC_6_678, I679=>output_MAC_6_679, I680=>output_MAC_6_680, I681=>output_MAC_6_681, I682=>output_MAC_6_682, I683=>output_MAC_6_683, I684=>output_MAC_6_684, I685=>output_MAC_6_685, I686=>output_MAC_6_686, I687=>output_MAC_6_687, I688=>output_MAC_6_688, I689=>output_MAC_6_689, I690=>output_MAC_6_690, I691=>output_MAC_6_691, I692=>output_MAC_6_692, I693=>output_MAC_6_693, I694=>output_MAC_6_694, I695=>output_MAC_6_695, I696=>output_MAC_6_696, I697=>output_MAC_6_697, I698=>output_MAC_6_698, I699=>output_MAC_6_699, I700=>output_MAC_6_700, I701=>output_MAC_6_701, I702=>output_MAC_6_702, I703=>output_MAC_6_703, I704=>output_MAC_6_704, I705=>output_MAC_6_705, I706=>output_MAC_6_706, I707=>output_MAC_6_707, I708=>output_MAC_6_708, I709=>output_MAC_6_709, I710=>output_MAC_6_710, I711=>output_MAC_6_711, I712=>output_MAC_6_712, I713=>output_MAC_6_713, I714=>output_MAC_6_714, I715=>output_MAC_6_715, I716=>output_MAC_6_716, I717=>output_MAC_6_717, I718=>output_MAC_6_718, I719=>output_MAC_6_719, I720=>output_MAC_6_720, I721=>output_MAC_6_721, I722=>output_MAC_6_722, I723=>output_MAC_6_723, I724=>output_MAC_6_724, I725=>output_MAC_6_725, I726=>output_MAC_6_726, I727=>output_MAC_6_727, I728=>output_MAC_6_728, I729=>output_MAC_6_729, I730=>output_MAC_6_730, I731=>output_MAC_6_731, I732=>output_MAC_6_732, I733=>output_MAC_6_733, I734=>output_MAC_6_734, I735=>output_MAC_6_735, I736=>output_MAC_6_736, I737=>output_MAC_6_737, I738=>output_MAC_6_738, I739=>output_MAC_6_739, I740=>output_MAC_6_740, I741=>output_MAC_6_741, I742=>output_MAC_6_742, I743=>output_MAC_6_743, I744=>output_MAC_6_744, I745=>output_MAC_6_745, I746=>output_MAC_6_746, I747=>output_MAC_6_747, I748=>output_MAC_6_748, I749=>output_MAC_6_749, I750=>output_MAC_6_750, I751=>output_MAC_6_751, I752=>output_MAC_6_752, I753=>output_MAC_6_753, I754=>output_MAC_6_754, I755=>output_MAC_6_755, I756=>output_MAC_6_756, I757=>output_MAC_6_757, I758=>output_MAC_6_758, I759=>output_MAC_6_759, I760=>output_MAC_6_760, I761=>output_MAC_6_761, I762=>output_MAC_6_762, I763=>output_MAC_6_763, I764=>output_MAC_6_764, I765=>output_MAC_6_765, I766=>output_MAC_6_766, I767=>output_MAC_6_767, 
		SEL_mux=>SEL_mux, O=>output_row_6);

	mux_row_7: mux_768to1_nbit GENERIC MAP(N=>32)
		PORT MAP(I0=>output_MAC_7_0, I1=>output_MAC_7_1, I2=>output_MAC_7_2, I3=>output_MAC_7_3, I4=>output_MAC_7_4, I5=>output_MAC_7_5, I6=>output_MAC_7_6, I7=>output_MAC_7_7, I8=>output_MAC_7_8, I9=>output_MAC_7_9, I10=>output_MAC_7_10, I11=>output_MAC_7_11, I12=>output_MAC_7_12, I13=>output_MAC_7_13, I14=>output_MAC_7_14, I15=>output_MAC_7_15, I16=>output_MAC_7_16, I17=>output_MAC_7_17, I18=>output_MAC_7_18, I19=>output_MAC_7_19, I20=>output_MAC_7_20, I21=>output_MAC_7_21, I22=>output_MAC_7_22, I23=>output_MAC_7_23, I24=>output_MAC_7_24, I25=>output_MAC_7_25, I26=>output_MAC_7_26, I27=>output_MAC_7_27, I28=>output_MAC_7_28, I29=>output_MAC_7_29, I30=>output_MAC_7_30, I31=>output_MAC_7_31, I32=>output_MAC_7_32, I33=>output_MAC_7_33, I34=>output_MAC_7_34, I35=>output_MAC_7_35, I36=>output_MAC_7_36, I37=>output_MAC_7_37, I38=>output_MAC_7_38, I39=>output_MAC_7_39, I40=>output_MAC_7_40, I41=>output_MAC_7_41, I42=>output_MAC_7_42, I43=>output_MAC_7_43, I44=>output_MAC_7_44, I45=>output_MAC_7_45, I46=>output_MAC_7_46, I47=>output_MAC_7_47, I48=>output_MAC_7_48, I49=>output_MAC_7_49, I50=>output_MAC_7_50, I51=>output_MAC_7_51, I52=>output_MAC_7_52, I53=>output_MAC_7_53, I54=>output_MAC_7_54, I55=>output_MAC_7_55, I56=>output_MAC_7_56, I57=>output_MAC_7_57, I58=>output_MAC_7_58, I59=>output_MAC_7_59, I60=>output_MAC_7_60, I61=>output_MAC_7_61, I62=>output_MAC_7_62, I63=>output_MAC_7_63, I64=>output_MAC_7_64, I65=>output_MAC_7_65, I66=>output_MAC_7_66, I67=>output_MAC_7_67, I68=>output_MAC_7_68, I69=>output_MAC_7_69, I70=>output_MAC_7_70, I71=>output_MAC_7_71, I72=>output_MAC_7_72, I73=>output_MAC_7_73, I74=>output_MAC_7_74, I75=>output_MAC_7_75, I76=>output_MAC_7_76, I77=>output_MAC_7_77, I78=>output_MAC_7_78, I79=>output_MAC_7_79, I80=>output_MAC_7_80, I81=>output_MAC_7_81, I82=>output_MAC_7_82, I83=>output_MAC_7_83, I84=>output_MAC_7_84, I85=>output_MAC_7_85, I86=>output_MAC_7_86, I87=>output_MAC_7_87, I88=>output_MAC_7_88, I89=>output_MAC_7_89, I90=>output_MAC_7_90, I91=>output_MAC_7_91, I92=>output_MAC_7_92, I93=>output_MAC_7_93, I94=>output_MAC_7_94, I95=>output_MAC_7_95, I96=>output_MAC_7_96, I97=>output_MAC_7_97, I98=>output_MAC_7_98, I99=>output_MAC_7_99, I100=>output_MAC_7_100, I101=>output_MAC_7_101, I102=>output_MAC_7_102, I103=>output_MAC_7_103, I104=>output_MAC_7_104, I105=>output_MAC_7_105, I106=>output_MAC_7_106, I107=>output_MAC_7_107, I108=>output_MAC_7_108, I109=>output_MAC_7_109, I110=>output_MAC_7_110, I111=>output_MAC_7_111, I112=>output_MAC_7_112, I113=>output_MAC_7_113, I114=>output_MAC_7_114, I115=>output_MAC_7_115, I116=>output_MAC_7_116, I117=>output_MAC_7_117, I118=>output_MAC_7_118, I119=>output_MAC_7_119, I120=>output_MAC_7_120, I121=>output_MAC_7_121, I122=>output_MAC_7_122, I123=>output_MAC_7_123, I124=>output_MAC_7_124, I125=>output_MAC_7_125, I126=>output_MAC_7_126, I127=>output_MAC_7_127, I128=>output_MAC_7_128, I129=>output_MAC_7_129, I130=>output_MAC_7_130, I131=>output_MAC_7_131, I132=>output_MAC_7_132, I133=>output_MAC_7_133, I134=>output_MAC_7_134, I135=>output_MAC_7_135, I136=>output_MAC_7_136, I137=>output_MAC_7_137, I138=>output_MAC_7_138, I139=>output_MAC_7_139, I140=>output_MAC_7_140, I141=>output_MAC_7_141, I142=>output_MAC_7_142, I143=>output_MAC_7_143, I144=>output_MAC_7_144, I145=>output_MAC_7_145, I146=>output_MAC_7_146, I147=>output_MAC_7_147, I148=>output_MAC_7_148, I149=>output_MAC_7_149, I150=>output_MAC_7_150, I151=>output_MAC_7_151, I152=>output_MAC_7_152, I153=>output_MAC_7_153, I154=>output_MAC_7_154, I155=>output_MAC_7_155, I156=>output_MAC_7_156, I157=>output_MAC_7_157, I158=>output_MAC_7_158, I159=>output_MAC_7_159, I160=>output_MAC_7_160, I161=>output_MAC_7_161, I162=>output_MAC_7_162, I163=>output_MAC_7_163, I164=>output_MAC_7_164, I165=>output_MAC_7_165, I166=>output_MAC_7_166, I167=>output_MAC_7_167, I168=>output_MAC_7_168, I169=>output_MAC_7_169, I170=>output_MAC_7_170, I171=>output_MAC_7_171, I172=>output_MAC_7_172, I173=>output_MAC_7_173, I174=>output_MAC_7_174, I175=>output_MAC_7_175, I176=>output_MAC_7_176, I177=>output_MAC_7_177, I178=>output_MAC_7_178, I179=>output_MAC_7_179, I180=>output_MAC_7_180, I181=>output_MAC_7_181, I182=>output_MAC_7_182, I183=>output_MAC_7_183, I184=>output_MAC_7_184, I185=>output_MAC_7_185, I186=>output_MAC_7_186, I187=>output_MAC_7_187, I188=>output_MAC_7_188, I189=>output_MAC_7_189, I190=>output_MAC_7_190, I191=>output_MAC_7_191, I192=>output_MAC_7_192, I193=>output_MAC_7_193, I194=>output_MAC_7_194, I195=>output_MAC_7_195, I196=>output_MAC_7_196, I197=>output_MAC_7_197, I198=>output_MAC_7_198, I199=>output_MAC_7_199, I200=>output_MAC_7_200, I201=>output_MAC_7_201, I202=>output_MAC_7_202, I203=>output_MAC_7_203, I204=>output_MAC_7_204, I205=>output_MAC_7_205, I206=>output_MAC_7_206, I207=>output_MAC_7_207, I208=>output_MAC_7_208, I209=>output_MAC_7_209, I210=>output_MAC_7_210, I211=>output_MAC_7_211, I212=>output_MAC_7_212, I213=>output_MAC_7_213, I214=>output_MAC_7_214, I215=>output_MAC_7_215, I216=>output_MAC_7_216, I217=>output_MAC_7_217, I218=>output_MAC_7_218, I219=>output_MAC_7_219, I220=>output_MAC_7_220, I221=>output_MAC_7_221, I222=>output_MAC_7_222, I223=>output_MAC_7_223, I224=>output_MAC_7_224, I225=>output_MAC_7_225, I226=>output_MAC_7_226, I227=>output_MAC_7_227, I228=>output_MAC_7_228, I229=>output_MAC_7_229, I230=>output_MAC_7_230, I231=>output_MAC_7_231, I232=>output_MAC_7_232, I233=>output_MAC_7_233, I234=>output_MAC_7_234, I235=>output_MAC_7_235, I236=>output_MAC_7_236, I237=>output_MAC_7_237, I238=>output_MAC_7_238, I239=>output_MAC_7_239, I240=>output_MAC_7_240, I241=>output_MAC_7_241, I242=>output_MAC_7_242, I243=>output_MAC_7_243, I244=>output_MAC_7_244, I245=>output_MAC_7_245, I246=>output_MAC_7_246, I247=>output_MAC_7_247, I248=>output_MAC_7_248, I249=>output_MAC_7_249, I250=>output_MAC_7_250, I251=>output_MAC_7_251, I252=>output_MAC_7_252, I253=>output_MAC_7_253, I254=>output_MAC_7_254, I255=>output_MAC_7_255, I256=>output_MAC_7_256, I257=>output_MAC_7_257, I258=>output_MAC_7_258, I259=>output_MAC_7_259, I260=>output_MAC_7_260, I261=>output_MAC_7_261, I262=>output_MAC_7_262, I263=>output_MAC_7_263, I264=>output_MAC_7_264, I265=>output_MAC_7_265, I266=>output_MAC_7_266, I267=>output_MAC_7_267, I268=>output_MAC_7_268, I269=>output_MAC_7_269, I270=>output_MAC_7_270, I271=>output_MAC_7_271, I272=>output_MAC_7_272, I273=>output_MAC_7_273, I274=>output_MAC_7_274, I275=>output_MAC_7_275, I276=>output_MAC_7_276, I277=>output_MAC_7_277, I278=>output_MAC_7_278, I279=>output_MAC_7_279, I280=>output_MAC_7_280, I281=>output_MAC_7_281, I282=>output_MAC_7_282, I283=>output_MAC_7_283, I284=>output_MAC_7_284, I285=>output_MAC_7_285, I286=>output_MAC_7_286, I287=>output_MAC_7_287, I288=>output_MAC_7_288, I289=>output_MAC_7_289, I290=>output_MAC_7_290, I291=>output_MAC_7_291, I292=>output_MAC_7_292, I293=>output_MAC_7_293, I294=>output_MAC_7_294, I295=>output_MAC_7_295, I296=>output_MAC_7_296, I297=>output_MAC_7_297, I298=>output_MAC_7_298, I299=>output_MAC_7_299, I300=>output_MAC_7_300, I301=>output_MAC_7_301, I302=>output_MAC_7_302, I303=>output_MAC_7_303, I304=>output_MAC_7_304, I305=>output_MAC_7_305, I306=>output_MAC_7_306, I307=>output_MAC_7_307, I308=>output_MAC_7_308, I309=>output_MAC_7_309, I310=>output_MAC_7_310, I311=>output_MAC_7_311, I312=>output_MAC_7_312, I313=>output_MAC_7_313, I314=>output_MAC_7_314, I315=>output_MAC_7_315, I316=>output_MAC_7_316, I317=>output_MAC_7_317, I318=>output_MAC_7_318, I319=>output_MAC_7_319, I320=>output_MAC_7_320, I321=>output_MAC_7_321, I322=>output_MAC_7_322, I323=>output_MAC_7_323, I324=>output_MAC_7_324, I325=>output_MAC_7_325, I326=>output_MAC_7_326, I327=>output_MAC_7_327, I328=>output_MAC_7_328, I329=>output_MAC_7_329, I330=>output_MAC_7_330, I331=>output_MAC_7_331, I332=>output_MAC_7_332, I333=>output_MAC_7_333, I334=>output_MAC_7_334, I335=>output_MAC_7_335, I336=>output_MAC_7_336, I337=>output_MAC_7_337, I338=>output_MAC_7_338, I339=>output_MAC_7_339, I340=>output_MAC_7_340, I341=>output_MAC_7_341, I342=>output_MAC_7_342, I343=>output_MAC_7_343, I344=>output_MAC_7_344, I345=>output_MAC_7_345, I346=>output_MAC_7_346, I347=>output_MAC_7_347, I348=>output_MAC_7_348, I349=>output_MAC_7_349, I350=>output_MAC_7_350, I351=>output_MAC_7_351, I352=>output_MAC_7_352, I353=>output_MAC_7_353, I354=>output_MAC_7_354, I355=>output_MAC_7_355, I356=>output_MAC_7_356, I357=>output_MAC_7_357, I358=>output_MAC_7_358, I359=>output_MAC_7_359, I360=>output_MAC_7_360, I361=>output_MAC_7_361, I362=>output_MAC_7_362, I363=>output_MAC_7_363, I364=>output_MAC_7_364, I365=>output_MAC_7_365, I366=>output_MAC_7_366, I367=>output_MAC_7_367, I368=>output_MAC_7_368, I369=>output_MAC_7_369, I370=>output_MAC_7_370, I371=>output_MAC_7_371, I372=>output_MAC_7_372, I373=>output_MAC_7_373, I374=>output_MAC_7_374, I375=>output_MAC_7_375, I376=>output_MAC_7_376, I377=>output_MAC_7_377, I378=>output_MAC_7_378, I379=>output_MAC_7_379, I380=>output_MAC_7_380, I381=>output_MAC_7_381, I382=>output_MAC_7_382, I383=>output_MAC_7_383, I384=>output_MAC_7_384, I385=>output_MAC_7_385, I386=>output_MAC_7_386, I387=>output_MAC_7_387, I388=>output_MAC_7_388, I389=>output_MAC_7_389, I390=>output_MAC_7_390, I391=>output_MAC_7_391, I392=>output_MAC_7_392, I393=>output_MAC_7_393, I394=>output_MAC_7_394, I395=>output_MAC_7_395, I396=>output_MAC_7_396, I397=>output_MAC_7_397, I398=>output_MAC_7_398, I399=>output_MAC_7_399, I400=>output_MAC_7_400, I401=>output_MAC_7_401, I402=>output_MAC_7_402, I403=>output_MAC_7_403, I404=>output_MAC_7_404, I405=>output_MAC_7_405, I406=>output_MAC_7_406, I407=>output_MAC_7_407, I408=>output_MAC_7_408, I409=>output_MAC_7_409, I410=>output_MAC_7_410, I411=>output_MAC_7_411, I412=>output_MAC_7_412, I413=>output_MAC_7_413, I414=>output_MAC_7_414, I415=>output_MAC_7_415, I416=>output_MAC_7_416, I417=>output_MAC_7_417, I418=>output_MAC_7_418, I419=>output_MAC_7_419, I420=>output_MAC_7_420, I421=>output_MAC_7_421, I422=>output_MAC_7_422, I423=>output_MAC_7_423, I424=>output_MAC_7_424, I425=>output_MAC_7_425, I426=>output_MAC_7_426, I427=>output_MAC_7_427, I428=>output_MAC_7_428, I429=>output_MAC_7_429, I430=>output_MAC_7_430, I431=>output_MAC_7_431, I432=>output_MAC_7_432, I433=>output_MAC_7_433, I434=>output_MAC_7_434, I435=>output_MAC_7_435, I436=>output_MAC_7_436, I437=>output_MAC_7_437, I438=>output_MAC_7_438, I439=>output_MAC_7_439, I440=>output_MAC_7_440, I441=>output_MAC_7_441, I442=>output_MAC_7_442, I443=>output_MAC_7_443, I444=>output_MAC_7_444, I445=>output_MAC_7_445, I446=>output_MAC_7_446, I447=>output_MAC_7_447, I448=>output_MAC_7_448, I449=>output_MAC_7_449, I450=>output_MAC_7_450, I451=>output_MAC_7_451, I452=>output_MAC_7_452, I453=>output_MAC_7_453, I454=>output_MAC_7_454, I455=>output_MAC_7_455, I456=>output_MAC_7_456, I457=>output_MAC_7_457, I458=>output_MAC_7_458, I459=>output_MAC_7_459, I460=>output_MAC_7_460, I461=>output_MAC_7_461, I462=>output_MAC_7_462, I463=>output_MAC_7_463, I464=>output_MAC_7_464, I465=>output_MAC_7_465, I466=>output_MAC_7_466, I467=>output_MAC_7_467, I468=>output_MAC_7_468, I469=>output_MAC_7_469, I470=>output_MAC_7_470, I471=>output_MAC_7_471, I472=>output_MAC_7_472, I473=>output_MAC_7_473, I474=>output_MAC_7_474, I475=>output_MAC_7_475, I476=>output_MAC_7_476, I477=>output_MAC_7_477, I478=>output_MAC_7_478, I479=>output_MAC_7_479, I480=>output_MAC_7_480, I481=>output_MAC_7_481, I482=>output_MAC_7_482, I483=>output_MAC_7_483, I484=>output_MAC_7_484, I485=>output_MAC_7_485, I486=>output_MAC_7_486, I487=>output_MAC_7_487, I488=>output_MAC_7_488, I489=>output_MAC_7_489, I490=>output_MAC_7_490, I491=>output_MAC_7_491, I492=>output_MAC_7_492, I493=>output_MAC_7_493, I494=>output_MAC_7_494, I495=>output_MAC_7_495, I496=>output_MAC_7_496, I497=>output_MAC_7_497, I498=>output_MAC_7_498, I499=>output_MAC_7_499, I500=>output_MAC_7_500, I501=>output_MAC_7_501, I502=>output_MAC_7_502, I503=>output_MAC_7_503, I504=>output_MAC_7_504, I505=>output_MAC_7_505, I506=>output_MAC_7_506, I507=>output_MAC_7_507, I508=>output_MAC_7_508, I509=>output_MAC_7_509, I510=>output_MAC_7_510, I511=>output_MAC_7_511, I512=>output_MAC_7_512, I513=>output_MAC_7_513, I514=>output_MAC_7_514, I515=>output_MAC_7_515, I516=>output_MAC_7_516, I517=>output_MAC_7_517, I518=>output_MAC_7_518, I519=>output_MAC_7_519, I520=>output_MAC_7_520, I521=>output_MAC_7_521, I522=>output_MAC_7_522, I523=>output_MAC_7_523, I524=>output_MAC_7_524, I525=>output_MAC_7_525, I526=>output_MAC_7_526, I527=>output_MAC_7_527, I528=>output_MAC_7_528, I529=>output_MAC_7_529, I530=>output_MAC_7_530, I531=>output_MAC_7_531, I532=>output_MAC_7_532, I533=>output_MAC_7_533, I534=>output_MAC_7_534, I535=>output_MAC_7_535, I536=>output_MAC_7_536, I537=>output_MAC_7_537, I538=>output_MAC_7_538, I539=>output_MAC_7_539, I540=>output_MAC_7_540, I541=>output_MAC_7_541, I542=>output_MAC_7_542, I543=>output_MAC_7_543, I544=>output_MAC_7_544, I545=>output_MAC_7_545, I546=>output_MAC_7_546, I547=>output_MAC_7_547, I548=>output_MAC_7_548, I549=>output_MAC_7_549, I550=>output_MAC_7_550, I551=>output_MAC_7_551, I552=>output_MAC_7_552, I553=>output_MAC_7_553, I554=>output_MAC_7_554, I555=>output_MAC_7_555, I556=>output_MAC_7_556, I557=>output_MAC_7_557, I558=>output_MAC_7_558, I559=>output_MAC_7_559, I560=>output_MAC_7_560, I561=>output_MAC_7_561, I562=>output_MAC_7_562, I563=>output_MAC_7_563, I564=>output_MAC_7_564, I565=>output_MAC_7_565, I566=>output_MAC_7_566, I567=>output_MAC_7_567, I568=>output_MAC_7_568, I569=>output_MAC_7_569, I570=>output_MAC_7_570, I571=>output_MAC_7_571, I572=>output_MAC_7_572, I573=>output_MAC_7_573, I574=>output_MAC_7_574, I575=>output_MAC_7_575, I576=>output_MAC_7_576, I577=>output_MAC_7_577, I578=>output_MAC_7_578, I579=>output_MAC_7_579, I580=>output_MAC_7_580, I581=>output_MAC_7_581, I582=>output_MAC_7_582, I583=>output_MAC_7_583, I584=>output_MAC_7_584, I585=>output_MAC_7_585, I586=>output_MAC_7_586, I587=>output_MAC_7_587, I588=>output_MAC_7_588, I589=>output_MAC_7_589, I590=>output_MAC_7_590, I591=>output_MAC_7_591, I592=>output_MAC_7_592, I593=>output_MAC_7_593, I594=>output_MAC_7_594, I595=>output_MAC_7_595, I596=>output_MAC_7_596, I597=>output_MAC_7_597, I598=>output_MAC_7_598, I599=>output_MAC_7_599, I600=>output_MAC_7_600, I601=>output_MAC_7_601, I602=>output_MAC_7_602, I603=>output_MAC_7_603, I604=>output_MAC_7_604, I605=>output_MAC_7_605, I606=>output_MAC_7_606, I607=>output_MAC_7_607, I608=>output_MAC_7_608, I609=>output_MAC_7_609, I610=>output_MAC_7_610, I611=>output_MAC_7_611, I612=>output_MAC_7_612, I613=>output_MAC_7_613, I614=>output_MAC_7_614, I615=>output_MAC_7_615, I616=>output_MAC_7_616, I617=>output_MAC_7_617, I618=>output_MAC_7_618, I619=>output_MAC_7_619, I620=>output_MAC_7_620, I621=>output_MAC_7_621, I622=>output_MAC_7_622, I623=>output_MAC_7_623, I624=>output_MAC_7_624, I625=>output_MAC_7_625, I626=>output_MAC_7_626, I627=>output_MAC_7_627, I628=>output_MAC_7_628, I629=>output_MAC_7_629, I630=>output_MAC_7_630, I631=>output_MAC_7_631, I632=>output_MAC_7_632, I633=>output_MAC_7_633, I634=>output_MAC_7_634, I635=>output_MAC_7_635, I636=>output_MAC_7_636, I637=>output_MAC_7_637, I638=>output_MAC_7_638, I639=>output_MAC_7_639, I640=>output_MAC_7_640, I641=>output_MAC_7_641, I642=>output_MAC_7_642, I643=>output_MAC_7_643, I644=>output_MAC_7_644, I645=>output_MAC_7_645, I646=>output_MAC_7_646, I647=>output_MAC_7_647, I648=>output_MAC_7_648, I649=>output_MAC_7_649, I650=>output_MAC_7_650, I651=>output_MAC_7_651, I652=>output_MAC_7_652, I653=>output_MAC_7_653, I654=>output_MAC_7_654, I655=>output_MAC_7_655, I656=>output_MAC_7_656, I657=>output_MAC_7_657, I658=>output_MAC_7_658, I659=>output_MAC_7_659, I660=>output_MAC_7_660, I661=>output_MAC_7_661, I662=>output_MAC_7_662, I663=>output_MAC_7_663, I664=>output_MAC_7_664, I665=>output_MAC_7_665, I666=>output_MAC_7_666, I667=>output_MAC_7_667, I668=>output_MAC_7_668, I669=>output_MAC_7_669, I670=>output_MAC_7_670, I671=>output_MAC_7_671, I672=>output_MAC_7_672, I673=>output_MAC_7_673, I674=>output_MAC_7_674, I675=>output_MAC_7_675, I676=>output_MAC_7_676, I677=>output_MAC_7_677, I678=>output_MAC_7_678, I679=>output_MAC_7_679, I680=>output_MAC_7_680, I681=>output_MAC_7_681, I682=>output_MAC_7_682, I683=>output_MAC_7_683, I684=>output_MAC_7_684, I685=>output_MAC_7_685, I686=>output_MAC_7_686, I687=>output_MAC_7_687, I688=>output_MAC_7_688, I689=>output_MAC_7_689, I690=>output_MAC_7_690, I691=>output_MAC_7_691, I692=>output_MAC_7_692, I693=>output_MAC_7_693, I694=>output_MAC_7_694, I695=>output_MAC_7_695, I696=>output_MAC_7_696, I697=>output_MAC_7_697, I698=>output_MAC_7_698, I699=>output_MAC_7_699, I700=>output_MAC_7_700, I701=>output_MAC_7_701, I702=>output_MAC_7_702, I703=>output_MAC_7_703, I704=>output_MAC_7_704, I705=>output_MAC_7_705, I706=>output_MAC_7_706, I707=>output_MAC_7_707, I708=>output_MAC_7_708, I709=>output_MAC_7_709, I710=>output_MAC_7_710, I711=>output_MAC_7_711, I712=>output_MAC_7_712, I713=>output_MAC_7_713, I714=>output_MAC_7_714, I715=>output_MAC_7_715, I716=>output_MAC_7_716, I717=>output_MAC_7_717, I718=>output_MAC_7_718, I719=>output_MAC_7_719, I720=>output_MAC_7_720, I721=>output_MAC_7_721, I722=>output_MAC_7_722, I723=>output_MAC_7_723, I724=>output_MAC_7_724, I725=>output_MAC_7_725, I726=>output_MAC_7_726, I727=>output_MAC_7_727, I728=>output_MAC_7_728, I729=>output_MAC_7_729, I730=>output_MAC_7_730, I731=>output_MAC_7_731, I732=>output_MAC_7_732, I733=>output_MAC_7_733, I734=>output_MAC_7_734, I735=>output_MAC_7_735, I736=>output_MAC_7_736, I737=>output_MAC_7_737, I738=>output_MAC_7_738, I739=>output_MAC_7_739, I740=>output_MAC_7_740, I741=>output_MAC_7_741, I742=>output_MAC_7_742, I743=>output_MAC_7_743, I744=>output_MAC_7_744, I745=>output_MAC_7_745, I746=>output_MAC_7_746, I747=>output_MAC_7_747, I748=>output_MAC_7_748, I749=>output_MAC_7_749, I750=>output_MAC_7_750, I751=>output_MAC_7_751, I752=>output_MAC_7_752, I753=>output_MAC_7_753, I754=>output_MAC_7_754, I755=>output_MAC_7_755, I756=>output_MAC_7_756, I757=>output_MAC_7_757, I758=>output_MAC_7_758, I759=>output_MAC_7_759, I760=>output_MAC_7_760, I761=>output_MAC_7_761, I762=>output_MAC_7_762, I763=>output_MAC_7_763, I764=>output_MAC_7_764, I765=>output_MAC_7_765, I766=>output_MAC_7_766, I767=>output_MAC_7_767, 
		SEL_mux=>SEL_mux, O=>output_row_7);


END behaviour;
